`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
D4j/ZvDlHH94W8+IJJbNPNXw9DmbJ0DFQqMp4WCxLo5qYzlDh7JWGs6yUUAdYPinbQ5v+f5jiZTZ
brp/kQyCNA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ndn8E8xYHccAX1+h/PuCGO09+WGamaUuTVsd8ob5bZBAgfj+wJS4buY6QgRSPkseI5tEjsLD5puB
988qwrfhhKESUoFl9yltwUtimd/sTAXU2WYKhQLEbeKvpBu39BTfXcEvLHplwONKXSFXN5ISH8Yk
SF9BM8Ula6noDPZAj7w=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XcXCPujxnxCyW90p5vBzeeraL7UcZpkRDUxGQbHOqtu/RkwBmTzWVtxgrzDg5JQIfNCk3j/Ir++m
D+Cm3cnjbceLRuVhF18NnkBjMvptHiwIyvdrTwhM3bbgccjUo/mXFjBPIOJctj+6kXD4hHJ7VzaI
h/JN+dwDzHjmtCDZzJ35NqPlrDrGHCN20W2pVnFqPXsNiwgOsCc72INB2yhO/xO5ajx6+yFMG6sY
LWCGLKL22wgJpdBiCZ/VxHWC6/Ay2lyfdmanHsIEQebGFmZpAmyrXpz6RxvG/Cud2ROTqutXkdwP
zReVR5t8T+nLd/GYRWhaTJ2kRsR/45yyKeT1jA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iyX9kBDU3o69yfSEqzSVamX1SVHKkjCVnXIwSOZ4UIgOoY6U1A1LEngp/YeceyG5cv+1utANZ23v
O5LWGf5tI2s9LyGaIjZ+sH7bHJZJaxMCoVke4gqtnofmcZE4PUUtqUHuZSrECWtFCS09VsH1+/19
EmHAJelN2YgDZLPptMY85j2zcT/fighjD3guUxdo3ZV2gUg1lcs1GbMgWghpdtT8eaf9DjUoBTSi
Ks0EQ0V9A24j8gL+k0/k7QIIpGvoK11X0jX4tFtSEophfBtQsEwKAhjjjZkp0xu2IXZN42KvgZLl
+P7gdrq4Ag3C6XJkRlJZJoypExhoDXADWtn7/Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sLjiN3E8+QLmHvk/t8+ljZWP49DrIBUTu1rmFpi/39NtC+bd0ihWkvptD5yKXIJWHAnj3pg7oTkx
wFcxIxGBVQziWV4X0Cy14L8AcNbfEpaUkcT2NRvYcTTe/igaLuQnD94f2kO122KfnbFzpPKXwgAp
qchh/EzggUV3ZvcBQuE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KlgvJ7nPoi6sNtTRWHdQeuWpzpzcdfnnVsEProzv0ZLVGjE4Huq/NcgICukVqgJEig/EltDssAFq
56bAlN7c4RkfjpwYF8rqBXH2/lt8Chbx797X/92SI/+nKffm5jdeEbZcNl1P62uVyLg+o7iEfpx8
lhdrQthrFvGlDCRTtbLEszl9OScFE54DvwrFle/2dlqL/qe+BcYFxueYCLweFEgLfXNUcTXVRr65
43k+osB1nV4lmWR7saLaFZ29cy1S7ikHcd9UXms/YvoEF8GGfmgcenmBPRQVKoCF15hCb/0HlR/I
eJWggCCa/nMGG9e9kToQhyWb6UshfeaWRGE2vQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PObFMgHuR7YzErHa0a2JXKTwbvGNoXpcB7tIVUzxyLGBZ8cJOMZlHK0ZnVzflfPcMwIb6EcLuE3F
Z9d4JWwpj8mJmyyU8Hqay9EMqH7UI3192wpiWOE6cJSjeTDzpwwg7wZDR4PPG+in4llvTfajo6oP
f4psWtDHzh9524YRzbgqrBkGo7yAOcJOJVziJWuuT2C/n/zl+azMb8sLIxSBL15u2/40pTLd8dL3
e6SqrnzY9JkUaj7p5VVc/danJ3zQJHhzE2Jj9aaGZR7yfX555EMxGaoTryvMpgTdDPePWb0hF9Ud
d2+atfCb1zUYjFS6odJETRRSPw4eOfZHTaeo/w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hOAgf4riFQqBBRwkLjpncD4vJLT3cULn8tK4LJCv1JVoSutwpzcWlmp7wzsD+LDz6VB1ugnXY+LU
xnyNmEzybWzkhXQaMc9ntL6EFf9+GK6tJrk2qVTVUM/JIUrsUO9LRJ/2ImUyD3bkALjgoIpXzrQx
98CMqi8XBf50ePane6UF+gLq7FLQTAtNK8lwSYb/KloeUxO5hox8DwMO6dP2255653L+Qyn08iLP
Oo6lQNxPpV3917Rh1Cg31uCfcbCkASkIT5aKlfVhhyRTefCoyRGzq3kgGqHrP4qgyylsVynlKh0K
aHMIVpHCH+SLXCFE3o4Dw62Izmwpo2UvLXSHNw==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SFXCXUmkNxG6cho5IN/jlAJ6rv7Q18PpVCuJlc1gcldaeLYITP69W70c+wznx7K6fqXVa1dc6f9Q
io5we006bznvtLyJv/CoIkraa6AxPihDwAvCv7/MVxL3jKkdYYWOBD2gKHOx6Y2jWKP5RcQFJUnC
Oowpb/NpxcCCyv3ETx5fNUDfxhtyov7hmt+YgkbD2WbTCYfrERIFW9T+f58TDtflC9otYGO8ILBP
YFzICoSuUpkggzbNKe0KRxTbUo1G8XDfqQxhpHytIjtCLmVj4ywLFAuh462lXvIJpextssnUC0Sb
r6zWwVuFIbSN7KI2BPsKsKKz//nHHm9JG/Rwag==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 566368)
`protect data_block
VkBFTCl1YgABFBOOoaUrVtPsLQMvVyYTnkdSl1gqKu0CgthEH0rxT4EkVnY5eZ3q5DFxtHkNz1YV
WUvxgG1mtaMoi57empT7mstZgxP57c+NsVswJAA0ZcpCScmLf5EX3ZdF6sBT0cVu4pDbS4IfLo6P
UPWI0RvpZNqoIknGsmL9BfWfQ37aQJ5T4o4gg6uHAtCut9MV9GZbNLUlD+AsWUzXnAaiCeTnxJPW
hBs4rHYIjA8yBaDVDETjeEV4MOnULBuvsSePvqcon8yOPABUCCDs9/ZvKFnRKxgR7it6hKWrsZmJ
fdMyJ94F+2yCA7cx0V1wsgHY7z7CbqEnYmt/x1FgAryl8bHjigCbA8DhxjQ+94wiZt6LYZO41FDN
aUJwsNBkZPkaL7vnbDjHrYZ2hWGI/P1GI7Q5RYVFVfLWqlpdVL7rSBv6R94rtpGH63NtfaZqhiJg
g/5OTsNK4b3iSMQhbU+V5Ct+p/BUwJthEzUgPajLV4QGBFw+hd/00hDc5WYNYNuID5JQXKGalqpa
YTA8W9NnhKp2V8DJkpUvrOoV8b6+7LvHL27R1qibDFbBk3ursaj81nJ41HQ7pd4al65wLUuUJn0x
MCox0rxtnE1ycTsxS4C+TSq4Lod60ASNDcnR6uYKQ+Ci5qPZeNHUs8fwzT5zD+268pBNrTLvFRny
Yle3f5EJGTOFINYW38tpbXgyz57WsQuOIzcR0Rhoe29aGogNhNs+jy8+AarlWmY1Sn2JpZzMdP4a
J30TNvTFs+eUWUN73MkCkyPhcFIiEdFlrMnYC2/PnV3lqWW3iBVA5LUXBWc0RC8zGkDnlwwhPVLu
y63FKj/xmP4D0nYif0ypbXyY5e8ERw3slrTn/QOsFqD1GNRNDU7VDLz7x+ChYeMGFBBRv1odByoA
kQ2XbxMRVnbJNuSjmi8QTEQOdos7ypn0Rd6SNCH8PBdvlzl9hhmiwbr88Tnn+dM3z9ZpvEXKCtne
gKxE3pYjWoZGAYrbbhiZqvkfBxMuLD7WSYAvBgoVSQcaMYGhW2/9dUiyvi5z4ttHMqf+gRsiMNiu
980oxjJryD342mD4dXS8AlCL0zTIRgHIindOfbIh3srL0ykK+i5eTrvRpD1Hf3WTtXTp1NKGFNtC
3ZsyrZuWL2yYOsX2+ygmjLIejKvneoNexyPYpYY7EpmrqXRM8ph4ygO+tqxdAunaBA0dz3Qvc55k
acS3YR43SbO/7Q4NaCn5vICaunMbwJFectRBt3th1TjsuujgJLV1b3HDa5r0gnH4Brnu451eFoEI
g2DPPzUQ92pXzpVgy/Ogrgyax5p5gSh5cFo9xG9VNhvSloG4rIc3e9+Ce5O/YyNkYFOI0SORzyY8
NkczztQcTTuhttDVWBQbPsAI7tNjve2+zgtKXVMD0m64Y+ZMiLH/0b1Q65obUgRaYTmzIFEeWeDn
JTIFKzZDtalJpv8yM5ASM9iGncyVd5WM7On4frz7KFLMczc4jX2uB942wfdYtZVTqrK6THtDEX9m
QXdH2a/DGscIcuB2Vs+XANLv+qlD4EwDnhGX1HcPFp5i/Tu2sulNeCyuBfszosKD0LIfdMEHtCYb
Mah4DHK1ZT3hMm7mySe4F0faLizBKspB0Vs0mDBY/UGbDz6t2hhjrS8aL4Qj3gCHW3EA58t5GDl0
FLSmxQbZ1xoK4yDNa9UHxxD7gWO2l89U9gdVtt0FKZENjP0Sl3SDDp2LqTb2vvNlXlZ6R4zn99Gb
6WSmXkYMPkoSF6Fa0uv/QKtP6+00blENqzLJ55S2zkSoPgDhFW52k99bTziFw6Sb0ZJ8Wm2YAQIq
l37oOo1uyZlbBI/wd1r3fy+dEXUOqtbvecCVh3sJEF8bmQHKYrT7ANKXVpfU92jO+NG8dNh4Cyta
TmBxUfHCRxMckeGaEpUe1P3eO6Px9tLJeMUwpPoJY1j3h1RtL5LI35tpM8qrCwdNTz1Z99k2EaPu
sWMOYwQYGwSLjC7puXSDQVzPWdi8u3Tn5TQ12SQvqkfJh0QOjJ2Rs1+WIAlLZj+kTIJe92w4feGX
DynIB/aoV2PymB2OO7MsB8FPutHdwToHrUGXVX5S2SoIBb4yRqXSOaACyi8wWcCQfIKbhI1MrraV
tWBfUOT2OALKhyHA4l5Tlw9zeqxSF8jCuuoamt14dP7yXTrgVZqxYPzYutfBQlVX/FhsZLm10e3x
a4j7YMg7ndWxovboYkfb2CG4UCDTbpMgIL464WnLgwdijP5s1T4HDChyy5a4tLWa0o0vL/VwPmFk
1MohtC13X3tkg9czvX3IfMRTR+zLhopC5pR/KjTQPK2F3CrNciAso5qM7yGHo7kOeDv8rWUFVnKC
T8C2Qrq9+1Z2hUzV6LwtwnPZ+CZ/SdTxw4IBsAs5eQHrzZLdXUYImbGJ2eJe3s/DAQ9dSv0XrSVc
lJvajFFxO3BCHn9Uz9OYNIqnxgYXiephzX4iFE2IwLG+vwmE+iFBXjypyUnahu7y76/6rxjWdEZJ
8vQzJt0VaLpzai502YyvaxDly4dtCVBXaiEGKezctoqoxm1a4ZdYzNB4XBZG5wwBXaEdSi5HLCwy
1ec0CjdJ/59F7ZW3xWf+6jLSgcbB0uACllVd3s4Jm8W8yLV5d9xaEK1Vs7ePdZ8YVX17i9b9WwuW
8dln/Hk8tDNCSuNHn5iJvB9fHwZ45rX0uhZ9Mp6Jd70F5QW9DsYverNnh8rPuiVLrI/kGrRTajV7
7lh9ThUZKC2B/ULlFAy+l9TqYFuQ7/pAI69fPiCwhJQB0fE6ubj7ET+ql4+bpiD8vZODV/8sMDWb
S85BmwW7slSZZUXskOtnpPSvzR7O5W9K0a/Cct5GLx8DeqDpr7NRKJxIH+QMyK7i1L090HX1hWBn
Oth7IgUuXnRWYz15occy4sMagAs8G0zVgAlI1qaJKSEHY4kakZIL15ocl8gqmfs7UH/XnIK3DtFR
qdluHrrP4BufbJtS8N1i6bbbG3Dh3ys39X5KWRnnh1qlI1Ev2WVmgR1FyK3mSam9JOAooW7R02kv
GkOa8n962DZP74qTAEWscCl19ivHmltERqbmmGbZkdUjX+wkKCiXfyUbA/4uktCuGbEkCc+TWIjq
k776CqUwaGaopQrpXWvZWbttvTZEFqlvhHcvCknP6JeCVel4M8W6Wh34Dg8MTw/RVABnfb/M581/
BOJXB4geJXW+Kl9twzOEE13G+YNtqlLJkbxWbdTbvGDVz4zlWyNMqoD6harvW2H/yU3/D2t0B9gx
qB+2uC5o7o244k0g9HRVfN0g4IqPMNHUBGnkdylJwUU9/iY7d8dLVM0E7FZou48c5NFeNsr6wl2U
OoanR7jrCAVm5ItWviAAJnMa97wwbDx93uu4vcFu8u/bQ8i1xaslgTXtt6YIqEB0XzifFR8vL2rP
maotb00IApVYly/qxa9ruM9P4279Diy5N2IUUycIZi3yn2JhbgpyU19sx8l5v4JPDTynW+byx4f3
qriDCR7msyRbQWeVVj0lgStyTFRVfSYy9Sn/lQwilW+AzhhEyE71jdLMFosDfPC4fNkH4EdChqqW
Y98+PsDB7vg9budQUaH7RSFfLoYv6yBz3Uh8lh9PmXDFrmXQ6mixjihWaZGNJVUUGDhcehbb1xhI
d51TnJqLGCQCDhw7QTRHh2ZdAHpneNh5ubFfAYB5RP9aAnz95TcWW2DOPpTDOlnJ5vBN3jchHXv+
eYKRy1rvcj7v1JHsXCv3vEVEJT1s1cPIeo+MDHRCh1u71jVvDzm0eDiicdcNVyM5m2xJHH68yNqU
+uoVcbLxzFSzM7ZW00U4JlEwLkSut6tGhUkKNaHOmoHcw2nM5aaDnUuHABYp0zv6mZwlU9GVY+/m
wJuhGmZa8auugNKKyJTe+H+Amujy3SmWEufMJbv/9ePkeYU4/TvVO0QH8acbBV1ob7Qon11mPFmH
qlQXxsoDOmC1iDOgutTIiHZRCLg+9mU7ZmHP+xR5TWuadLm5MdloVZ1C8VtIKPF68bekymjY7u5y
HEcCu6qV73SbBdc7jwpoimBh/pLXLaLczBOw6veLj5fQ/S7/juQ6wu/4wkIieDKsPlHTgeo+RxkI
KVwDM8MUXirKuehXMn34cIqh7ZAnKo3YaVfsouihyChZPyQozZfAt/E8Tc3zka7cw/rbAij4xF1+
WM9lWsFNmzZS9uSHsTZomrMoe2sP49ok7wN4o0LK2Yh8sqUQmEQJpBOpefGBgIgU7rCTiwlzvmZC
DHvugguAUnze3SHFvuI7uOg3DqGTNqED+qlRRUvgpEu1f0qAZgKAx9CiTuVL0iv5EFnbVse9pS0f
Sw9HboAFnFASqklxp3ho5lzaDkySywP552EADI1L+Q3gQoP/DbaENfizB7H8ECKUkU4438flgbVU
Pfz9CukAPRDf6gwuzxA61znP7kebrjIpzm9AxVrcYGs01RIOy9F06jzSYbJxT5GzP1QUL2UYD3gT
eettj590CniAcWFGL9bgfWNTPcQ7R7pczbCUM2xaXy8izBccbrqr4wLZ0In537rbXo4r6k6MaEx9
l0D0DcUjzU8yub8EYgeCMsvSk+2ancri/lpCsKh9Zug+/WDHLAyfKPrPe/hmtQhEvsMfFm3lIcyT
QHGX/9n3d2P+nN6rG4tKV5VD/Vd9nIRTM5U8fQHtYLWxghC0CrznWU93tG9sS0ZzRcUQOMpHmzfw
6sptGhJ88toC+uZ6QPvsb9cgQ0zLfnj1KvWF+pvxl0m0jgCGGkJJ8ExZ+t968DyV7DpJxtDv+sHw
EC+qvdNXy9YyW4cRkNpqhkMP8qd+pZDR2LCN0gXDC6Qon7wXftMaOHs0rh1mSFKhnTfXpt654OG6
ImQ2YEU3P4Dke3/Loz8brwmYygoumgCHxpo7xroVDh0oIV+uPJ0mxcDtovrnsHWMszacnfaPlSsS
gkRvsczdc954klzi2zaUM2y/EydtlFIxdDNL6Yd8EVzAieVyGy2TwsH/aKOZeCTaSzO/j5ZSkPze
Z8/u8g1lDa6ET0QexAfTUmKMCjRAH4ZT5idq340bOVdDwP/TFvyafRh9BZlrGws2MupgYalM9pXw
LczD9t1maWfRLJ6Q8grOF5+taQlLwgojAnWOiA1YZ+D7nnrxXC/kaf+HuS/xbwUdvKgQn19EHaNm
m7DTJW9igSMXfRobaO9q9koWOacn28/EqvvJHztBhA03zTrXQVOxvolJhhtSJNzS+FQ4xIRzp0Wc
Yw185ETNXwgLkEO1ApUW7zN/+19eUCVNFt1v+N4jswFTmNmrmoOWg7kRJxGS1Q+dwCcphcVmyNmh
8KtLENDew5i8FksgkS0wwfFj8CzC1ay+bvWrYoMXj5QDxavomZwB/y19Tt86ITbipaEC58L2RZLX
YKGC4GIPTuNNMApm7rn7scVNWbbLru2JHHgagPrUw/JQK85TcXxzMxAGcyw+1Sw9Yfe3pRjHeqfb
Akrh7sNb4el7AzEABrXM+NcKSPjdwIh89Ys4fd/BAofisvWzHILBgOiEpCI/dI5eNiRn5jh3oqhy
t4xO2Is9WE/pxCmcslqTPkiMJ3IYOzjkAkQKDikT/WQFj1YenVP09P+fx6FGNrao1gGICCtA56Jb
xSRgFse02X74iywbD73nOKWEYIinA7en+u2VeSizzbxwmHXaJzf6waH4sfNHVSORelzBjdFDFMaC
/Jd3JMg2e6GTHIDM2IfBMRBm4FKkd0zB20w4ZxECqeXkcAommUbnTmneI7VITJI05b0gNBWQhzwI
aTkOmNHSUm/Gy5SaQmcJS4wYzhd29jrZws0aQS29awyUZK6ocUkV8sZ11Ihh4OLUoJ+0rl9hUbh5
En8opW4gHuP66Zw4vCw7TTO3DebymxEeIh0hv5/J1Ol3NCN1izqZNKi7KOBU+BKfqPZJHoJlSD/0
zuslCMKc03HxWZnPfp06s90nBRR0amEgQT8mJO8ODOyTt3rKhVAH5UanhxDmZc0p7UPx2gJtVwJl
zzFUjyqOoUUYQjo0ZoOuNdOr45hn4vCa7/3F2U7GaxEETe7RCprPlzmoY/Zj/gRgHX/hucIYzvGj
4guMQYxre5CItNOl1p4zyFDgE5eQ5Ls4IUi82PhC7q8Uci2iHxkXjzgMhb3M/avL9J1gU+o9A+cD
L/mTr+If5eoq0xQe+TjSJ8PGJA8Ci7jQhx3DGQpaE3Q6QDcZiJYcqgrWf5xUkb+O0yD2r40iGGHY
EA/10vofwNUkKGkH7EO6EkYOlaYKvTLHzWOHqRvBxzjCl/D4DbWzkrDtx1BdPYJsJ20xkx4DqlNm
PItONPLsyk8wc5IQd+be6M5NpyZ3Y+DCWHof1m7PMYK6YsOSSRVIX8aFr8NFEp2Mkw/DSnBRSQQz
A0w7NzCJYFFe4Jka3zVHdcuXtPnJOVm5ifjqS/SQn2ryaBafXEBUhOXQ2svkKzsfAqdIzdr4zKcl
j3J5KNagkm8zABedt4YC9+UIWFNKEvE0lHmx1bIAyuSFSmcaroDlgXHPA5j7YyZi8q0z/0yVSZOc
mvclzPp6cmKbr5ltUJrVX8dP09YJ7vTco9B517QZPkbtXn08Ffkksht4hoXYIWcpT3dAe0qokDFd
K9TVmihVy7INOwTwLKY5W0G00LZfhDfuqN63nNtmZVkycJ0mgb3LJ5GZQT2azUB1BjdFaLhyT4KR
4PlhIKeZ3Bq+lMrbf0HIpSYa/q6f2RA60EqdWvHvJ0hGCbO5zkqo7kOKmaqbC4/vny+4dC2Wsf8z
vebQxllw+BngrWl9r/ic2xc2hqbhW5+HNPGyK6nznC58MYJEEuNKFRNXTbj1cN/iQtPa/4XMGllA
DR32P2bmnb9G+J53l61iZp6GEUpRzZlVPONslLtC0Vxbkrbdx/cORZCbRQRb6vgoSINaQ/INR4Uc
eUETadIuYKvZTEMPFtdzrxa8W/n+oGmEFxae+D6bBM1NXNP6QAOra6+in6mpHLMZ/Vl6iQZwW13Z
pC464UYoHPO1SGxjCdH1L9GhFanWQISahDtwntkfswG8D86yzhOsGrDJ2iwEVtlJVLBx0ee293L0
whKdMnQ9BRcwIkDHajtti/q1UVlK6FnxRhL7ZNQmbfYswPguFHE+3ep7sCiz6CrSTbVDgy/ZMO1w
qTtevWW6MHn3ozx7YERZPeCdCFcnrEhQCyZBVCBt6L6on3pIhPeSKd6ZRgTmQlX9alMwVT8d4UVf
cYlE6WTODrWI73zaOXzuB4RDa6dMIHqhQpUCIqnGicSDRjehUMV4dO9Mnpu2QuASW80fK5M/99y1
ocH6QgUcXS76YjFHGu8cRPsYIS8r3m2Ts/e/t6dBGhvTIVwhywfF78t3+SH88uFU36qd04aVia3g
lhBxVzFjqcEIYixgmvEK+ajtXtBwBOQeP0+MgYl4Ga5i04mhaZlDl+lFRXIMlcXjbFYfpF8OW9Qe
p9E58jDT1c+MQAfHuLSFOeBLh6mwvQFHXl5ycTpY4lDLEMpcnluM6vSSTPjkHn91UQk7N7NN8J3h
7cpG3A1HzTQn+moBgcUPMiPVpKpVN61DgE9beElBtYEfjWklfm2V6CDBvQBsUphUG/dupcyjlsOt
qT1+7neB82crvXI1+2bOtZy/B8Bgn90K18RTeIDpMhSJS8PB2LxSinJVjZYIpy0g73JkvDI5pgOM
XhWq1pHWN4F0jDbZZMSDzKcm30tjM8Fi5udgkOODfvyfJM/wZJQuXxAu1XK8jJNfxqfgvov5PFke
MdJUvEFu2Qs955uMBO1teSglAIIJDr8XtphYchOfcd5rDmWtSd9Qif/awA9LnatFjc8TYqrCCqoO
zCsnXhmftS48g3ZsSzZGEIDpcF4kIGGIA2Q+zINvBJomF+/tPuKs0qXk5zvn7Nv/GcOHqWnrxbYh
rC/UKL4EMw1bcJ5MyBanGJzvfhjhKrs3whUnvPIu+SdyCEo+LnjuigZ/tG4982rNZisTxS3jT5io
OYs9+5m6wceNwUbNf+1fB3Ri/q8a05UPGJw73pzyK6uAEOGeYn4vcgwi4286vojse/hXnL+XHz+C
g3CAn8XXMdN+i5oE7nzflFGnlWcZEapXatqlQIAS2Jr0V7UR5BpT6ryf0IQCLj+NJoYREtSBvJiC
5VpdHzS+Qu/kJ2qqZw0xxMed0O5p+yFedyt2JL0+lV4ZILDS8lL+mnoJLIJju3k0du2alnjwzvqt
Mkkqa208xDlpnPvzf+4SS/+WoACAWnzR3X6KsaiYt3KKKezAdaJ5Ap0qJitJWzIjdp1sWyGPShDg
bwlUTQu9py8rCiDNy6d0X7nYUSUpdDl26RVJv+6NkRd17sGvewhwoZ7TBYwfwDEl35v5NPrRMR0V
xn/qcJq/8OA4YtdJH5UzcKVTd6IbJc7xCNn2BNI+mIVmZKFBrRzpIF4oQBi22euysnGsPYroFjj/
rh7Wtovxo4MR5q10v8PVqRhIPXDlwKFQV1NHnmFbsQ4aHToYWBgetmemPKy0tsCDbT8c/MvuZRlT
4nNE66GDP6d8+ZnVVLk4m1+dHpK8d+Opfuo9mkSg24XibepH0NAYfY9qCDLXFpMyap/QQnhwbbd+
DW+YKZgnMyQ93YD7hTFTJ3MNPtuwx7F3IjHRausLcIHvnWRyc4xXGVUNt+VP9CVzpTc3jpJtz8vG
YyrArfcqu4/l+eXDV8pSsCxosE63z2hTF7ESQdDm88l3OU0WJR04xd4JeFIuGwSNKeYuboy0GMMD
FnXOJAQGAFVv8/YFCIj++GrSrvpeminbYdE5/XWmbKeN55VIdCJTFfqJwAX/VA61AIRdVh6l3vnM
wvZK2M6puNH3yQmw56QbTTSLDy7tbQa0ex0GqHcaB83GwmHr8cPfbINcc+QFTLkI1qMAGxbQWxyG
JvM0nVAad4YZ7ggzBYCqmzhmAattA74qODYSrVrE1z9En2QMguzDehJPJ/6d3xFIKNyyYW0L2mVW
7wyrwzvyMtTXdNebe9eMuy1Ecvc1eDvXv+Z4xdK9T9iObx3JfvQTlHnszB6rg1FNY6XzzseTprzI
hdO/TTzVlAejR9uiDeRopsi2R3llEAMZ9qV5/bixkPBNyZsyN6BhfcQpHtrx+Fi7I5+huW+WlEuf
TzVtofse4vEO5oIxEobunDptMSvsgksQVKUowTyr9QGITs3WqCaQkXie95Ap+wMf5OA8DqJiSn0z
+mUPfP2ViaZ5WZ820TliyofNYqMMprNXhduiJwpMcNjiMsTb8QTbTXy5LFSR31a03FghSyVSjY+r
ry3dnv0iHngETEzFIqe7ZL2aYxiJC4pCqTP0ZW4ZqfDdKndBD01I8UXehUYEF8L/rLWkx6PbjDxD
92xCnrN55l5awbmumMuAs5jF+5D2isbHyJtQGQNRsGv5sOTVnKfmfooHS6Eqw0/kJahf2i4UmTiv
fdL1Ln6qgsLwpEoWLnSxr7XLXMToAjyKl8GuZJk8VJHlJu4meocmentgUF4bgyWM3fsz+NXZy0ZJ
qKS/CJCIfp8KBQUuZAsLNaWAWRFUqD7arXLrjKAT7dcQR/v3yI07uZ1a2eJ5FBxoGPw7SHnILni0
9XT24D2gp+Y8+ypzAh+al8WC03nGW87346Npuxbapn0oZiEHrZqdqhmQ7bVt3JJGv4ggHUNgpvsk
Sy2tagT4P/OJlPC4vRX2ip4Agf6meNpRIpqF36igOuglZt8vwyO9NhcvzfHiXBD8kB/HdR+qVjAS
sBy0W5jNdvV0S/rbcGB6k+xPSRKtFETtcjgCVLIzZuQR4S6h08uB7KNw0CCJtY2LNy5AM0AGVE38
qjiamaBZZ3/6JKoXbkW+CjECiUBPCfELjFlE2wPxbW0ypwfEi3AHGBTQx6MAZop9297VZuhEPKUn
FAzKfuH5OVuPjDbm7gALcyIfaoYYvBH3adiGNI2LpaDSnEbfcm38PrfE0wmx5k/kHVi6RHgDEoY7
hEXwLdeqH9niCq2qZr4F9qT41Huc72OC3RsBEx7Z2A3WiodTEvIKbKJYDZHcNBCJLsmPGsCqDKIX
PWmqrcRnIkCzLFYRQ6JMbheCcYHCa/oSlzTGcjr1NqJAG0Brzr/SmwQodptNW0nuJrmxURU4kXf0
6qZkajiD+ZelBLrFRKIW9WPig1DCj6cpVa8bqjccCCujoo5GfTqwqDjyWyKD7wRznmm+9nay/Y3Q
QYbmCjsjxLUI2/Pw8SvQtigr6hQBlY0zO9EEFLsz7yqJ/ckSaxFLcd31gyupMSyLpDtYulIVP1eH
QwLIInREiYhNjKu8jz6/X1Yo3mO2EZLUihRpzZAIJNBFgyUZ8mpy8PG3XEI4cmt95NNoDdgWOwJv
sWRufgc0E94yx6G6yMJy2x9IS3ZYYDD5TVOdJOI57zPUKg3otAi2S/8K5kw4e6UtbRxzSmNeHxUN
KoRL2mCPZrS7TJRD2aj5BiRfK3C0Y3JGDaTq9fDagjZFkRSe5909bxyDVa50Yeg15vRAMWIYcYxC
50UcpN5sF10Ffimwmot9+ryYQVKKzcT9jigFgFsYfhgujkHjfeumHFG9eVafmBRuD4YNH9FnFG+N
C0htUwj22O/yTk7XB1g6j2jyCzkpB0qvVnNDhhQHh+UiQxrWdp/cwqYwTIzQnGMB5n+DtOyyyy7i
a7nONeXiQA3cOIEYhDTiYvAb3yGv4RGWepMhRl3/z2ilpVr6dH3goaBirHSwkM1fgoAo1HFx1iUq
stlyfTNrwYfupAtLw+aWwj31S+VxhmYyzuDJ0fo2HLFtwT0AI2GkQU3IxTK/66j0q4IoRtuZM7CB
w7mk//Z7rvWPhWee8c/BgEI5eoe3aI838bIb9QpiJirM9DLabGQyHoGzr441OEYd20/Q/Azrq6c2
Cs0OvCJ5bBgU1ND3HDJlz7tlFo80ijmMB7SUxFag5UvdwAP+P4Oi/7SrtMZX7+vfnXM07BmX1NiP
6JFOFSubNW7m+pzNiSTYSb01dJ3Gw2l366k8fRmcTVCd0D7qbcsngS1CYzKiYjUS3rMwaXBUg4Et
TlD4V3MUjrnaJD9JJDgjuDSFPHjEDDttIvwnDWkpKdNZYqGkBVfFk+PjFHGI6yTaX84PxhFWFx/D
IdkNdXIve4exPeG+1ZgspYw5Gajj9w237JuplPTKCbrjaY5bEZfPtjYsS9ppRMPBBrzMuIbdt0b5
M1HUOfcHhlhpyZDbCV1EHC/e/I1RCm9RDqP9QTRLP8pkPKF3Txgwe76Estm3pyIskKn7fam5mw4J
GLYvAzfGHJTUk2zjI7LBzmZPrPPbdxCjnAF7Q2bEYZTPCCE2186OgtjmouPGnijaqBzLofRl9KmH
AZmpLAcDFyEJAvSfSjrGmULFJBBVMKEJqP2D63bXC/C4NvhWFSe6GafarZ7yXAGxaW9e+Mj9yJh2
BKxsgLlejb3n51HYOOvV5gHX7Vk4zQ9lsuFuPPpY+drNb3K87dsPiQgw050zitvb/JH/ws8+/mHn
Fia7WV2tf7TaAQqb2p2lp7uMcyEau/NSC2GWM/WIKtLggbQahgliY94Xw+nMsRiCsERwVnDFH8Z8
xa9jo9yzLiRw4OAMdV7mhNMJxtJaxGf9HeXe1N6f8U677T5jSVOBokUvW/lu6xOg1YtMWeUCnF4U
CgR5kXXuSZKJnoqbsx7RTLV2X0va03RqDIaSPUL5H1zW3d1d3pb3X7AtRrF69005TZWLei+K75t7
7lkvAe6iCOFUIMi5zw+JhV9jZ4bEsirU+arVVI15A6WVqIRa3O4II3ZsPUzouC97P/S3QlacIxjr
BKn09+8WP36n4EKNZ8YDJM7VVt1EsnhGEDM26uIbtYPaYZXWcpiS+Pv05C5I/pKBY10Ah5pX3Wtk
vwIJh8FkTpfcaxYQehU2R8bw/OkLSkzKw8D/OTndqpfDVUCKQWLgfbKNt32V3ectjEGk+dx11iIa
H8vOqcGUEQvnYIoLYrTv10cKuC0rnlOQX4WUWdkO4fdvSEnCK7PLASuL3H00cg/SXZ8TYQHd1mS+
VNIMHU78qYaezvE43xQS0JfVfBgmk48IfcCdmPL0ISInf9fGgZi4Q4SsUMmK6b4aPz0hgolNpBM+
DDnh9O21KDB6ioxcCTOAy9PL7ViwNWtuy4jwC8mbViXmbfjwqGTIZQMnDojZJI1/kx1dlHSb21aP
SDumPw2W3x8hcGE+tjZsmK/GHaN0xRTSMHw8GworrZYh4oCUIplo3W4/8MSVkcbAWLp/r5v4ORmj
7FJdqxuKdW9UWw65QvadJgD0KzkmBGz2yeMxw5yOeXkUmCPYABe5vRmq2RL0qzk77/MqmaANJwQQ
gyTgKAqfwQ+nsOJJqc/m+gfw0Bf52VhOL7CW4kRqjRTGWPoXKZlgDfP5YXs7l3oGg1yeRT7hwXD7
TnkySdqFdhPSm2EZlupH68v2sDaLLx1ygaAzO+QnQHvd7anwJCKNY3pKTKvvhpns1jjQB01JPGEL
YajiZ8fpzE/tplSG107TmyZKpwrah7VFuu5XNx5DSUgsqyM2vg6tRbKY/cQPhj/i5fFrD4eg9bqp
Noix+eFfc13rE7cLVLFYKQE6JfpWy8cjirwNxL7jOn7HZ86mdWGk8XOXqhAatbvbsedYkotELdvs
/oxFSFG2H0g86Kcqit6QNuk6Hv2OweiZwy4RasgCkE2woI6DXg1NYOxYVsZb6YaSUts4arHc85IR
NwrS440w48mqXJmTK1JgfYDrEgyX7A8Bq8eq2gY+YlOwfaCr3rxS5bNVeJ9QBkq98j1eZ94iVxJ1
sC22VK2/BczMD/A/Wokm6ajlbfW8OkDYkOMX3VpMYd5yA8xUXjAXHVHpFc8W/x9LjLlOWoqxH51R
e77G2tl/Tvcu7K69T9TlOI++K1cchogp3I6z1QDqvgHJJgLMD5XFHIQ/utTkgj2NfjNy4sED0fuW
v3NSSYjsVQHJhpDT/ON0uHSZjJNTJfuyYjyMW4i3t8EYivc8psUUAVT/fkA4X4/rpTHT03TgVAkC
6TNSVGunWT1pHg3S+e/7//RPjT2HjzeWvOdFEorEbIZES379Zvs2tG4UCsfkvJfH/R2GYv/murz3
qhnd1sNX+T38SAViCgesnhJK8uYePMXeFLzpWC0IwJt5q/F4Epq6zpVeEkb8Yrqyxa8mMXSrSZFX
fGFPFMnmet3fTFg0C+h8l4eHvWlhYi6EA4n0rSnpCKHrCReP+RInBdnDbQA/uqy6Y+5jHFsQc1cd
f+JlWKMo16oXcpjVbZol5fi45WIBqi5ux1zK50cbdzK51uZtqxFSSixlWTe9JPHiAAubFq8Tfjop
3bS0ZkgSBZCoE4r5Potnv4I1ovHh4KZ4WmW/MbTVFu3Z9lFdc8Y9ZPKZ+rdFmGptRLFXyyqkCiDy
WQiVLfOAkQkTBSkhYkVlNruZuS6D9SvI8Yh+9b5NLQ2bSyfQYr7xgvTjRUyA6YXMcXLUgVulqOGU
HdL8eVWmaLtntHePBOz2aO42HKc+C4QkQ/zoMTVcKpEriGNP3MhjBWCqtGNRrJMsVq2xEEI4w3U4
u7Fi7ndQ31ceWVXIpdyV+4RgD8+g+CPR/kHuzFT08GJcTXc+7OKEqZNwiuh6f98Hb9a+hLRNM2YK
H4zeFEo2qpGpBzv57V6ynv5QAMfgq0UZbFymIjNqb4pPjCNXSgTFO4hTVrfQAcdguNntajr5h+OP
VUeL6bsD1LaLo045rs06tCNHJIDOvpNu30PfUU63xfT5bhWkG1smDX9fNuBt1mAPdTs7xBeyimhA
uuZYoidsEBlFEBNZNBgbALD/mPMim5eHZWtz7yyyv8xdMtBvq9LnRBxftSbwShNSRpZStT/YnhQo
qneMUJRMjTz3zbZxcLZbybX+UTo1y7i4tf/RIs6j1e482UM25vbHYy+VT1XmYj9X80Yjzf6eFsy4
IRZEGepmmFUhUfhU8KFMd/yJ77bf2XRkDURWd1StRaHLEP1KWzfM1qZF8JA97Sy3ZkC/PYbBoqUz
Tqtufparnoz0WR2m+dEXvf6k9cknpuLB6nQ2RjFkXQ2Wo+lqfr8lhwiuRehbtXTuD3dPNjMtmxZf
da4GVg3yX9xWthcNCQuUuDJ4OhybB5a1xAuof4dWtOJz5yVS7OtCtekrbn0mpyqa/hKQ4KSdOT9p
SGcCc6bFme01LE2Uxw3KqPTM79qh1v2zWL8lXsw8HZtfdqg+NJzaeD43q+C4LRwElykSgCYz/6F7
HfD9mD9kmr6dFZWcgSE/xbXdbjZfW/g6tjMGvAgXx7wU7jwFM3yLuv3z2m/KOT0Ae9ceO0J9dMCu
ksRs9qPWeaEZht0MIwb7tZHRRWB787qBfEr7u4PDEz2QHhpxCqSaOVA9Hn2Qplwf1JWlYS0GhM9G
K6+kOUMg1KzwhR6ryUWRTaBZBnzvufY4SEGyZSsNOhh6rpzeObxOyCugRBK6m5xENEruncXGdlSn
UajWffR0c7oUUqUuDF813glyiVyCLrHM2XYWhbQwEJZfMnes/v+IQCG9BTmWiSnE6bvWBTueq3I7
+g3lOYI5YjmiPT2vP/+HQ6sb4+nEaxE470Kbt0L+6K7zKD1dyPS2hKGo41PJYXRbSKEagONpUhkw
3e3Oy3GauMknPHKEILmXo47UFr76eOE2y+9s/PljzEAQKvj4SclTpfLq3lRwahvk9kfBp3ONsit0
m2NpD6ux07Hvm/w6NjerJo6wXeByzqyNqneHZ/xxjyxM3cduA6MyTVFfb+8929GHZ8iZ8R44anRP
VrjYW0tEU3BgwzJxjs/3QguRc3GDB/S11RsQvNELuvbNgLtprwyge7OunnU+xv9DAlM+SMfurin7
QQJq/jPb6byp8R/h9G1gUW4pBGj9cpYsxEAK5AawNWPs7sqEwAopju7gZlm6CHBuet0bIT3zbgaH
ANS/S5XXE5JA0rYZ2Q0emkCf+5Z1KKwg0duEVyZ54emUVhwJT60KDvfnOE53wLMiAy3lOJBYcHjp
U0G1OGtWtnTvS9ty4gza6OYW3TWgDLbhyoJIaKTW7xKYo0aNuE0F+1fzFMDezUgz++UVLbwBiViQ
egWGhM8bInMnG1JbDDns0qehP4XevjeE9PKnONlnp+kd9/gnxxVKuaMFVkGUR/Qr55G9NmAKoU7t
x1RRHgnOZPF3Vmpocn3AlfzH4DDmIjVNtsk1wBlddx35z1fqvgpkKjJ5v0RrEQPtaq0eQszQ+F7Z
h4MuBHjD0k1KN87TacC8JW1xHxqdLkhCtRt3uYXSgWVzzlwe7GynWC0MtLBkwhgqJM/0YzyVa1Ky
WxAgUaiY8YB33dF1WVOwZI0qeovS8oQGo7cszwgSktLDXfuMKSPzj5a0rPxsF473SGlsY2HBv2N3
6ovAFT3kdPOC7gOIFBIT3ixov9Z7z4TGcUBFsIczQPr2yNu3rnasUEarNAd50Ub9lqXDRYKKTt2s
XEwaWAaSUFmg1b0wmBO4cW7oLyMGv2Wv74t/I9GaJabiBpOjqg1ydWFXK7XpTdLEfkmUz9r/KVOX
8CmG9pgqwXTmaLMgki6vSwqr4HNVOPMz5bB+PbEl1GY2gPxQLQ1tIX+/O44rloUbk40dF+K1vV83
3z0hE1zbzBRRGfBPQ5zmgKooPs9Hx7DEElJUylNpU/Qnbq9le4M5LsQAO+r4tv+inh8TaaweUL3+
PRAeFId/O0aDvtnScKZBppdpah3etxb86ERKyxLfHJ8YAEiy0jKRpaf79OlfMav1xPwtVBENBnOF
2516BR30j6sgRZNlj6oZniOwuppZTB3Bswg/G5bWywT/bUT9bS6D1EyNRKMx4Vr3ImlYwBR46Zyu
IpCanq+DRyEySxMb9ETRniEFn7GnjnjuvzT19kkO6frn08+7ZxnhW/l0TLdc0ku7GFAaS4nnpni8
h4ppzR5OdwZKdZyMfIbE2zexpj8J1fVcKK7Z3DMuSKPXvxPAWphRsNyS+3wZMC5IEETMvfLhK2d6
ODur/yGVJUMfpr4N8+5MhghSjCfooLcyeoCqhpVSJ6DDL8XYT3ZBy5dNfPdmtD+gR2wXw42Ndcde
AvyZF+bdrthl2hhTGRuuln06/+xWrTPV9aZAXHm8lCzvlUNr+2eJWfhG1c6zxF/LsQYRjZpSzeY+
9d7Q7jj60Lr8CfyjibLXf2nDR6tAYkVFe06hVeKJ/jDJvOmlYBrtE5YXmF/eMq62kCkLcEm7XRFp
fcH8YAtUePRPlqSc4Sydg5GhOd8ph0pSj4uRJwh22xX3ULlrmKxciyZP3rx2RteZWC8gG6DpVp6G
ioorjAdo4iBJvnbTjxUSNv8GRsHrE0GyHQV3hL052nH9cN9S7cBXIxgkOodPfaAEGp8sjYJ0Pmnn
JqkG6PHlNwlnJw+L20tiYIML7EmMNIRWpMDLJBfjziPkJuyzqZahZmu3fmibhn7AOENc6I8KFvKc
br8j6MD8PxDD0rQxp5Mw0oe9NoegKi3rQxqqjcQLRLpG21gq6iQZAc1opgdotHN3+DIw+Vo7IqCT
kjqILYZv9Gze9Of/D0AFY18wMs6tlz+xxahg+hJoFXWJAxlKp+J5VmpSVTQ0SjJw+tzOzYlTXQ5g
IQWK1LXCNcM/cBnoDna5wrXd2yqgzLL4ZCQNf3Ed+cf7oYh6C3NReDlSQ6cUmM0VdHaGpRBnvOZb
oB8XAw3RivT0iPca3AIgldzi1JJAudFvLwObanSn8jBCK6LX/joUPWYGURzw/50DJwQBUevEi/rs
wScuXYjsuKaLzgdOR8sag0lbfDwrvLQV/to1mUB9buehGaITHyFl3Xbcwg3ccujKg5xum5BY7lrE
Nd0/Mta44Z3DhQlcYDFLLpClHfAkGY/6f90QzWvXJI21CmpFuIDCYyrpug1nTNazj9SIdf8Doyzi
yySsNYxcC/uSgxiL0LH7qldZhKBMSxIN7HZlu/pFAk4RnMUrkZjd4x5omMIGYfo6wFGhmVmkZxSR
YHL8QzUjUs3fQlIWhdr9MrafCGTMFC4rDFajsdBHw109IQAMMUvejG6m4j9Hhu/F+KSY4mTLZS3b
P4xqZVeZcsdoYIGkqJId+oYu77mBwRgmSx3vNyoCg22+JAOPgjvAQM7ASUStk0Lrr2KUNUKxJ3Ah
DKIDvBfJuxMn7cCn1z3yddilHLJmkuODmIQMpjZ9v9JoPd8SQMk56y6xY3AbovMyoT5cTpYL2HhK
eDmdJMLW4LUUGQl6b/BqkPUVfRnaqwTJtYXpRAC/N0sqaKWTzXkkmupVvqq/zkizNzhADVVqI+Gw
4olqLQkLc+rab/8+wjnOBgVzwjCb+x1HMyD6powpigl/2+PQp2yN9vEbULjnrkYDE9PecO92CL6B
DbkTpmjQHn+Dtmwnv9ZET/B7M3uJXD9bLnEkU/5N+mh0f+y/Kq0JsK/JC+L1fFmdS5V2sTX7hra1
9GXbKESpmT+CapwxNQne3oh6FV75lhs8h/etNIn1D2Kc3+P7Xa+xVmfM6/nW+Bht7qKtdDpVeM1S
TQivVGdpP7YiCNou0+pv3Q1rkRKyKrXUMh3NlhouXwtwexiUg6s3kNWSOympXXaed+V+wxroM1Ve
Gib2itPrxD+/W4x6YYhZZXgtrk0Tw+5GXOd26LXYoAsxo1X4Sth72d1KZf8Ze5grATyQnDo8l1or
XMNyTbh+RT5QZvle3EQ9Q2Pfdk57WrxyT2C3kOccMed3JT37eNGgPuuorvNkEzwAY5pKRzEfaneR
eN/JTdGokj+DRV7FzcY2TsNZe3/85FHXPgs/xtK0XwusbwyYL+2v6RoYPoPWEtQwsyuLlfe0DOyF
o1qq7iLPGv8TGas61ZCAoMQR+adrm0UVTy4nHJ+CIprL1HKxqB9LuKKYMKHQKE48HZaTJNbcCvEf
5bfdkV5stFKolLWM37vwoZHIZcBtEeASgAdRAUg8AZ7+aPKtB+0OukVzrpLYZPfNi6f4Cy7D9mVm
2Kng6EuV09qrdk6n/k5TvE3oVfV/HWlLYNhOALOw6yNfhTq9pWMfQ8iF/wlcCPyX8nmeQDSI0o4V
5EOjtJt/uCm5+10y0IjUqITnanx4wED/98Gp4p6UKI6M3ax6FW1FBc2hNBv6g+NCCW2vt4O3FEbZ
VNLzAEtC9Wmmt30QrpXZaWv79z3SojAQa9T1Yyy2zM3LiVsu5xqSwnrG/FnyLs2yWH+3Kw1DLKNJ
Z59ReSP00KjSe63mC5FXgtblaESFFjBT/M+LFPiIU0sORUuF92DfOguMOJ/SpTY40M9Hz5JFH/dZ
YTTjE2fpVlejHY6qdvFHGTTK3/J6wiq80KDJWCeqOxMaL3sMyBF+FbbEnljl5G/mJwINLpgplRBU
mnWf0/mk3ufwHtli6U23/jiZc8gw3CTuDZBGqG9YoU+RKfwy5oI6nr0VDOF+pj85chPP+IVhUB0N
s1QoabPIdoc0ClF8eAxtnBG9YROLRyWgN2OT1+FQoLV9OaLf3uIQwSmiVgESzdfPnPCa1NO8jCyi
gYyEef5beWBB9kHZZdlJKmPP61oPszqyXrnbrf7EQMLlGRU5zcAXtl6qG3JzIg/SG6thElx2wJ4y
zWWngDRfb+UDQNgvoF5cSO5uinGzlt0N4IiToneJRZbjdlz1iO7xfL+gjGgxJQy2JhqeslnYtKND
Ht5PQUrwJc2KL2tP/2WZYGfAMcyQ0+HbKpVb90v6lUjAPNEgGKlIsTN+29grO8vkw1U/CJ3u3yto
B2Ai53T6VI3y2iMQ2nltp9RMev7f3sfTDkmAW0P/BgBvuROm5FLpwLArAxSp/khrQO1zChzWOEMt
I0pjh1DgQzHmu2EFG0+XDkVOQTQQ317rEu1tODGGUuTydi7PkZIDSPLuqhFNQWDGLNaIEW/82kj/
DMFReeBGjnp2B2+QXo46FDs8m0Ig57qNZ5hyK0D9nhGDiHAi0Y06fPPo4uK3B4uzLRbSPe9sXT5e
A5b/JZgZPtFnAXY7nzb1pM2mx2tGakwrlN18xX1zOUn12bTwlz4WDbJQB07GaXPoXqOfoi7n4tGS
5tt5bEJdGbeCXQlEGlW06BIhNViChMILq8Rp6wtCdmwFFhV7jiKKvRnE4w4fBdsPt7j7w5MLDrnP
YBpQPVMlxYuvHJrw8lhiFr9g2y8SDpqBE4xBu1L43cbddRs6rxfTWSzvAQHvRLBU2U5ifttm6e7k
2JldAwGVtLjXXWevcZhylcDEvgYT9Gn+zWMh1yWWA8DkUtLS8rSQV1EVmP6WGD7DlSFj0L19XnrE
gbmERRz8Y8ZU1gk1Yw5PnHMh2HDcY9BuRC7yeA7foVQyN2F7HCSD812tzeS7eOxC/aEY9M9OEi1g
QkIKwa56v6TkD/rMrERYmQRbh5vKg6UJBDpQ2YhOLtCZkEzuSFvxlp/E04H4JUC66jnN8SFdcAAh
R+UfohgEDOmCnRp1aqA678knM7tQAOmL0kfev8l/GfD/EkOHM67j92eZ5gtNrAyfKWjmft0wZeTx
bOE6TlSnnTFNktDA1x8n9c9aXWg80/KYfhvQ3BosJvPCfbEoWDx96438yjrhnZFov3++FyesY/AJ
Ymj5l20SGWH8SXmCLZ14cQ5ZMDmbR34nsoDiTyMhsMch9eL+Ba1OC7dEcM/1wSA7h9tTVMtfXmnw
M9fYWdjcTpWOd5p6KXNIH/tPgctZbDYEoIdgH00q0D9+xg1bbgMmi19Xwz2cEdGMKjq/WX1dYvOn
GHA+SFE51d7YvX58+XOyXBEkJXKCKuW7TYVOApSx+Ic2fnsA2QeB/Zdt+QIQLzpovKVgFAOPgxoZ
H5lpxqMkNjaSPsGuB5dpTG9W8HLLyeTKDdnz8CC0qAG2cEdCrG9Jc0eI6oQ63YGxQ3VQJbNi7sD1
/XyaB3X87JUO0E0vXzNU0ZUWWdOQsRKML677dvYMDU5qx3KxpcWFoYivyf5a3vdWLd7sdEkJwmqj
2wBi1QWTb820+sfTxHrTFlBLVETWRJTTlpIdFfQ9XvY/RVcGeUnEBSPiJP2nMKrlA4Xiwdh4Bfcm
2aImkfJcTaLlU32i6e7pxdETqWfBofg9QwiO1LrzWd8/lpOcg8JcWT5GOeRux8mObf6LnWXnFncF
L1tbAk2kTdItoeVTdGhhoozp2fEfQnb6mi8xJdGsBcQMLvoqBB3FFsWBMUSNdeEMttNdDPRWnEHf
OulIuY61cZVQT7dM4A5v2xUCONOqIETaWCZoNYERuBUx+JWbLwOwd4yNaRCSlU5qy7S7tnzxeelL
ZHT2Me2AsE4MsYsdfkV88U0Y4zAyCJI1qOTMg35FdeOh0fdvgW1uiakopIujEJAnOhHUTwN0s3hd
PYJrMACSjLJcgnra0zKqP4YD/Ap3UainahopnIZg1j8FN16Q09FFRMdRtWsVUP0u8NhX01H0FXJG
ccN1uZ95UEH3EcAf06H40FeflVeIRbEXWq2J+UIp2rRgtnnn9VjR4qJgl/uW7TNRwdFlA1wB7dyC
rc99htr0Bfm0GKyZ7AqwSAZ3nB1jIDfE9h5KyExio8bvX8qX8Ah7cdj6WNkzvFoZH4xW+gpbE4j6
4NdRSiTuQoVbtt23AjlOd+KaybwvCPoFyVexsAvpqmoLDnU29OTvN0yQFdMmTMiWYsfxZBe2475W
uGJyr6nXw+HtsvMfETEsvaZKL2sv9cXbObcvdbpUsLUP/iiLaHkhYLSK3/5tRNUU98niep/tIENt
roe1JxoL8jtTm3qUkT6qkGeE95E/vfecCdEHOreWO53/IxxPI8/3nJYD1vsWixOEheg7f5WOT5ff
TqSk8QSOP4cmZlUtO+ktABiXasW1WexfDFouOmYfCADWLHRsxK0YHFAg1f/7eUQexx3GJcXqLI1A
nGP6dj3nBY5EzT/p2++dwtarBMx2Od4OLzG2y2IcUouoEiNdsIV8M0hNIEva1hWfT+GpBvR98yuT
FBBmZDjzNuqOm4dv6rOLL2AaUE8nns8X5kjYbqX6E/U1cQc/Wr6/jjRth0ZAb9njU+qFtjSRl1EI
uyh5/ogfSxhItlCudRH0Ad+pv/8hsvaY4gFuCxpkVs2VhDqDbv03c+wdtxoUrQYSZyN+xqVTCZq8
ODyuqtWGGEfvSJynacliVS6ExkQsGEMkaLc/YEaBJR/LlzkoKms6NaW8laFJjuQA2+nSMw7gHSu4
sGYqe/4uVAP3qqJywzNynMC8p7t1iWQFOHONgWxRlxLwCuhu/C6Dm5Lcc03HG4A+OTGjB4522cmk
IbjilfsHQJz/b2Tu7ycLg5BdIpJpaDRgwaZvOR+Q2qo8D/QTBu6EUHbyx5a1Me+0rnvM1kqRQra3
EHDTcodHeGiPtGbKSnSzMG5s2IXfYO/IEHEjsJvUeZL/KbMTw4SQc3sqpWQKq5mL0Ac0wANasOnQ
kKzqgWE40AK2oDhL2HOQsCfHkgEY0+Up2yrcSfLzWpZB66knJ8kue0Urkw/72yrT0wYs9/TNQ0Ff
Jo6W27BY0W5xBmHBOo+DBkVuCDOA6FP7PZKhtAjn2N8AHtMkCBZQUDLQR4xirjFvEQVbZDzdorzQ
Ak6khJp/KwXkL3DIUbbRmXx8dM6Uy9bB8jWosLr66D//VmFCjcB4FfLErT1iLbZmKGCE7vbv9HbG
HjmEceUCZ1pOONBUiUUGGnkC9wuYcnCNynHAKc7MXghbbtyYHfe/ax03gDz8CZGAitXHWuSHJBYq
dkBk5r1mnqVz66QcJgdu0dqLdm6ASdTSDsMHDOwKZsSMSSbDEuyHhhCGsHA+Aw/B49Pl+aTtBZZa
2MWy3WC7wiHAvjI4T+hmNKJUSwskNw372MvE5rAPkWqShgMUzW/27XcYh2JL0WOcUli7rjdIzg1d
Zjzm3F+TsJK4KvzslEk3Urwrl3UuJtY+eEMFmi5/6eQrdgTXS7DeloVhPrl3OBIvfnPYkacruq7/
L1TBlLr4uNoFviNCx2lxSfM8j5G3G/HCtDKriN9oeb7pu+cZtLhN62vkRa+dtJlWUVpf8qVSPQYI
175f3FOfMNe7dHHE1mOx868srh3R+eYyMxNdczDGi5M5RDWGctWNVXychKkPfcteEfMZ12RQM/+H
sdxFd5OHEMmH7w64YjSGsQH7i0sMfuWOz2GndP7q+uEsxa4NJs38uv0tins+ysKGW3VI26bCNJx0
sTpbHFvvWK3VFpHsyJGMCtzVUB1PIXSVtk4MGpcTKXnY0Yaw2AtYb4rGhWjq4MgYL378PvTWRBdP
ud+zoKCvKWXd2o9Z1uYcch/K9hHIYIsmgCOAuANmi2+0ImGPGV0V0zstw+kLlEFAyUb1nCTqGuMT
u8ir4QrpkdQpDXbFroDh2Fj0z/PNyTfGS24m0NqD2w2TgAaYYTI4FKN5lEwPZxlfkzTyVdC6QmKF
SqKIsg3zOSszJ68QwOEYDNUsEwFpamVpFgmvdbmVCfOltfLY8laP2BHLIPnKLspIkF0iCssrwcGd
5cYEWV8hxC+tdlSZRQ5QbYi50jmj7MsK9ugX+PznmZ628XRk3JIbR93ItDKjYWFs50dukKLmphSe
4NAYF1s/TosGiryWFPyaipIiUDU5ekCbERLMLLgXSVPPxrcISinORCnHh2iadwazYstzEyH/s7LC
NIjlyoYeFH2myBc2wYQjGD4ATvcAaHwb2JPp/d+vizJYPoY9al+qD+Rnhs7zxucHI02iOIkpmLFm
buiOAE999YitMMHxZKQsBTbzOebPi5TtOqXUQHBW9OuGBx1/5pC32NBgW5gHdTjietRSfIzn/EmP
+JLPsFgMkkm0HIH/UNrTXmL4S/NyPBO3GdOwwt1axKfkFmf9BSSWxK1ISDsqSZYOMbJIsBXdW793
Zsge6AgoQSGzb+J+rPsXGw2pvoAJNT1IvW3qGIw5vt2l6lK0jfPcqSm9oAQpdZxhJsjvx3VpqbCJ
XoPaMORthUWrvv/g8mrtNJxuvrQ3qLh0p+kVzURmMt0TR5N7d85ar1+yzv+8yRX1OQvisJ9uxWC5
geaB/0d52/ZXtFhmUkUf08B70+kM84SXd6QqArTFVG6pGiFobfR/eE9UHEJVjyLQAMmjLLmSHxcl
c5IN6szBFtGs+dgfUZesVXQycGLJ4uGcMYmuJmP284SMsycBPSas9IAkVxZc9zH1ztbBOAqGqXJJ
yxbyW2KJJhEkci+i9w9M88bwsndVJaO5bDuVucti8dYwTg8SYewFvfZw6ec2Uywn3hgQEQ5UEZWo
Rl7LsD36zCTf153Fch0LjVo/XOGaBSrN+/62FOv2wCOV0ZGsSFx1ZT2+OccItTp3Lc5OxUyZsn1I
t6Pj0M6ErAGOZbFZUma+7sYZG+1cm4Tq+fgRomr9a0E06DOwDTzjmWitmHw4LPnuAki0+wmH3JVo
vbTyHHpct04r5wUXl7smOQeQU6xrkpOGstwOSjh4C3iI4MGf49FQjq/mG1Qg866JFfVdRcmpOhoU
7RFUQlla9iQpi6BRW0hx9l6NTdHFeMxe+sJHS2Bpxtlbejt2c/Yp4+L4BG3KNILN20C/ZTwnLtrM
cbs+oDSJ0NiVCDzXuTi0ZdlLtWGpAp6KWzW4uzEDOA+HY+Nlngs0x866UUCz41w1rpapl5hsaqLm
wUM5+960fzze3D4ViaTQaK0LZG72fBhRjpOpEwhi7ITF/V08K4wBzF5vlmK6BLLTUuKYKINYCU06
QrBpzb5MKykIkPP151lZ13D3/b4bot1OfzFErzCQU/MTXANiY3D4DgN1lxFlXpOPRg2/txJz7Z9l
enRb4GoMzwunEVJfcxMak0Bg8EJgfS/fPwR3RhnwVBEGM7W6CiAZ5Q004kIh+mvkj8OnuD16XzTA
p331ujES7q8bvd4nWm1FaCWt1uXLt2ydQr+JNwF7xH5thFyG++p3JyN7wuvNSdsRoYhm3c9bqLsa
CpSWFNlIze3xJn1M/dOwYRwTaILrEsjH3xuIPtHR/1o5Zgl8xfIzhOYvsz0/NlXFmkwTc0pklQwD
8H/GhaYZHZsrmpysjQQpPaoo5RzKDeWdwgGLZB2NODL/woRNM7AB2jPF7JGP/tESfrI2f4j2W/Xj
R0kJ0klCLRA3jjgTpNFEMr8U5d2mY7GVOrpNZJ4wkx/EOuCdKQbbtmZZT5qigYHXfmxQ/g+Ssv05
9LgSEE7CrwTitXPqViY3iL0wreS5FEOjqCmCwnVtueij542JNqTG7UyNTua1p0heg7Ik21g64BTz
dy5+d3a4EJ1Z9wPCLX01ad86LT12fdUn/1XVp1gLP6UdSPpZGSJA6o+qB8Q+n8zEzkKUoRHWLndP
qgi++UdLLOckeIi7puTL3O4xLyD8nFqXDq68WPh+b8x+KqaNg++ZoC0Ii6ts0HOvmYieXfC0nrCf
8RZawcHmHWhHbxWEGbEJRSTAFBFUdlJe4DlkeUAIpQewJdzt2R4YbewVTmqipmBiutsq/kC7CJYZ
n6V+Ts9en15KZT9Co0de23oAe0xNg5XSM43x9K5nSvVRICacvL/vdw4gsJkQzw2zJibpq6iaLnvt
TfZOs9ZgnK4FK7kh7h6qDVlb39dgUzyKhGKrGOnslMwHP2AhIt0tSJFhpkF6nTC5xDXjF/IntHtL
lB6VTL0L0bdIinv3OXxkY4fX84OD1gjKrm87XY4hjhFBuuWzeITAet8P4KA3XOAxXb1hyTdaasYi
7lkpP5xq+gJFURHCiy+anb3wtS6dv5bO9XykDFfH4eR7uZj/gYE+GiJSPfrIgK2TvvxHh9julzaG
pkhUj7ORnFLjV4YwHuC4Tzx4r6/ZRJp8TZ/O4BpFT7XNQILXp4iiTuSvJ8OZW2yw02dQSY3jjJH6
CK2m3+jEhYBb3Y+cLnb5hp1G+Um2TqLN2HdJTgWpxw68JWbozVFaS1Atqq21t6yI7uFYUgkuLsvb
Jmaad40jEAuZ+LzioQD5IZc0GXNk7NVvpGQrLAY1oMiwG2I4pia0gbI9JM1Fd99IWKfPADFaXN7h
TOynJ7CLxXyL1FXnMz6XndPg8eyk7xygA+G57JP0MBeJ36x/Rd+9HEGBfJPz71XVCG0Iar9qDPXf
Lup31EVaQMFrOHUfTK3ldrJktdfE4M8vw3yRkKyH6yLjBEFmOG9AhePPugHcbohXhZ6Q5oQLZBr1
02asVyHyeDTBPXuAYfCRq81JPBNKufSC8EFh1QCMLo/QSwDOwg6l3gal1RfNhaOrbRTUisBjm1AL
MTDx7ATmz7hEMfsWSGrsoZiscIMmrv32g5AgQJciM9HkxbyUSxtWIL8UMZBBWr12hZAylC+A06JT
PLaukfAWhH3zIm8TTEaWSCW4gcN/ovkk5aOGgVHzaY3WLzZ6kXTxQpKO/3DdCCnlIzihV9+GXrSh
DFRbltGJ1g3oA3GPMrwM1BE7REnAAzEC0iAMGCKXLaHyy64YuGNH2LLHigxdGUdYH6uwJo1KAo0l
7EqzE1+jC6A+MSTKh1/v2b5h+GEAGlHAMUsbzmm2t3F8GeTjjV/f7GQ46C3MIUonvrU+2mqJq2qS
B1L+T7Pfn31mWcDOQO/A5IPND8/WWgCjNAzGyEK9+yUH6Ufmo84G8Ol3WAOMkWpk4wUgCmAhOvsM
FKjk6FC50ZKGG4dlco8wqUhVEvaASMQAs3jzhFWhwDk+XQE90UMbE4ZYjBRdPCYzYpsWWj8iz5qr
m9tFS2sThejpcigcWs0le6SVTZO2stUg0lU9ExdQing5dOpp/rar6jLziug5U2iUDIqta+b1cOVt
oD7I4FxRAajRqXd9aEcDYAtEgogxg5lFW9ZN0aTbfooAk4K1M0R4QoHzocp5MBA0MR4g64wCvjZA
1cNzkRH3LmvPpc9E3pay7lOfnL8Dho6zmzBcS421r2XZmCZq49USLzeE6MifQlXqMtUWSGhhH2YO
C8DR4/GPiPA30K0PTlGdwZPUH4rq51AGAHmoWtq6O06+fRvM68ia5g1I8bRW+02EN42CuJcK+8dL
oBC5QqG+E5XcqFIn/bB9UtTyhLIoKR6KcmmMRR9r90qUpYA+QzywxGYfDj4iOgzTx5jXJ3XjKbT9
Wc0r9VOjhMplqz4sr0g9e8p9eoYdNNeETna7Mij5jnZ5EruxgiePXBeQ3933+O0MOD3qux0appZQ
MHpB5KT+I1MRQSlhVUlw5Fsl3kpFpXw2g5qffq+47Hicxz1BOGNidNjH4PCpW5rftK6Ns3+a0qOc
ZaldXFDVyoR+lYmu1tL6M0CSqmjyWAVFm9Hua7JZDdO4I4HpvLcA8ByFYnxjRHdyGqrTQGD/+8Kb
jDghxHYLGpguotzXJSMLxrfDHJpODHn0++js0o+OusLXjLGMcTrSLQgVHKtUjuBmIZm8juJBD/eS
1d+7r6HEFfbxSwd//SEjFdiDzdmbO6+3U76lYpfDZjXGkyqvb2R/vCoZbhPouKnb/t4mL64tGZh+
u+GizBE6JAfaeX1mCQS6izXTo4oqBqHpZWxezydubAn9MkMJe+axQm7P4gKyMI3lmVU3Zc4Cpe0b
gHAQoitI/Pw87us0ofMg76GES6IGg/CkbgYTKXE5K9C8BYcui8FJX0c0u9ttJfqCaDCvv8E3FWV9
SqKzgy2hQC9bglPuvwz5jC/0WugMTF7UmJAjznVCxMqyZXiSwfgDOkgbcGOAzmNq0yRhPygK6tqK
XpJi0vrH1XR62gm2fZJEV3Obcsc/oQ98493j7zZFJ2sHSg9VvA+vlCCREuuo+BBphrGnY7/+tbZP
jt8ylDQsT9W62KHZAgZwq8Ou9xDz/BrQQOf0Jk3tZHEfYTWCFLHIRlKiCr96e4tRWHyhGdWM3yxt
YYUz3ETBE7ets/v+fTuutyw2stiU3dmPud6hRbOLua+PXITzM0rpd8ke0s5TRFYc+I1RwauIxrm1
M3g9QClbz2844qi/TS/B55mOgFy0X7zaC1apu4YG2LLENZJNl43wBGiQ2eWxaoP2eFZHzc1aXjN0
ziK0Ng+fRgRBWdS7dinMRA7c5zoZKADQzbjgsw8RmXYC6OtJm1RSC+CLFQRvlQPRivo3rwUGQsIl
hYScnaskhmHVZ/lCo1W3vOt6ZrLB3GiqB7rtuaMfGXOpodBodNat+9IQeiHIFr5IsFoZBzkhzwKS
QK5BgAWgrfLUA2xHepjOdN6x3Ka304y/oWgBXGqN9Vwkaxq4rD8u74xPIwdq658zQqHbzcyu93R4
nLHUSaDrZkvil68nUAH6LAQsUrKz1AnUEpA9HfZlSglrXic2MreWWzCXWdAduP3ZbeeLAZ95kRH9
SgxOpSSK0BPLb+p7nmiWC7X0uPXYHhX6IJjbSab8eNwspQH4Gb80niBvA5uZT4ALdd8V78pIX/Y8
MRdmQ/oldTvax17ZnaD8Ven8Lg2LRvCIgza8BWmQeyvCEt2pCUnHrM8CL1pzK8ZUDO/KU8zDlRvl
ckcySzzP+ryjh1kSjZa1/wXPaxOLa2O0G20RjmVfz+b0aV+FGpwm61DEZoy5O4NhSYZNX0F2YTfx
mh/7LunD04owH5m98XFHmEIyg5QcOL6rCEWUb8miMEwz7aKCt7e3UjFrG3Cq/s1NvbYyYzMhiw79
4zLwuda69j8UhqLIr7z2I/dzJCbPqT/QANdbLAKVGd3+SGfSk2PHhwP68VrHNzGnyDDUr2ZN+PoF
uN9CTmqLVNv4puRixRagUTu8B1FykDBsHhNN0TM090eTfPR2Nylzg+ni9jif/7R4KU2t9dtZ7QSF
vL4eAZgWqI16Viorb7ggMmDxbrMlgxZLHvry0zisDghiJYvV/UHSQffzv3wxDO55X+KnOZxpcvqt
lSe+1PUYmbzgoTskB5TVK0tas5ig/TwCCDQXPmXRCV03KydFoZfcB+k+L6X4KZ3YzVyOswok3M8F
RGwX1/iqtkXF2jFAPYOTLUghXXEu5qh2EUfb29bkzPtXEsBo+ij5N/bzaZXheCyS3vf9VLyhmZ85
NHgHHp6zLCtMutsXLZam+UGThXNl8a2cf+IKZTtfE9gQ9sEmM2jJY/Bu2SqePgAQdhPglqFZ4r+U
vWpIBl6h9Hx2VSnc12grWqzvFiq2tqUxoiy8kOanUPobdMCYo0LPBe4yVz1HyhOR6M4PNSzFWLUB
CgImJR1TlOjZZeREb6ci/4Aw9SkqIr/6T35H36S/TkdTbwBX3wckIX9YX43ThoaK8TqyJ3bMEZmQ
QFtafmItlntLMThpsyuyB63Gfh7+YBI7H/jYd4qVrUkjPBhjB42qD5TI0cxI3cs3zc9+Z2QFRVQJ
ws7Pbvni+vmX3+QPihIhrjbmDQBDKaY/vb3VSn9aQ+yuiZm/GgOg9o4bAlV8SZ82or+J7mTue6mn
57XLfgX5m0WkfhRDximylJTBfiKKbJb+xfleCmwKP9wIY2x9aRuFA0BJP7dZe+j3if3xiD0APczo
vbiH5voAvteTeY5n3NxFVJ2vloN63fAahdTqZDdVprIvoDh2iaUMYMTc8YWzQaz5axS9zKvBmhre
iwYl0IbPpXxNw4zxnRvrMwNXXhtg+4xcXBljJa4OALH4+Ta9VPa+AJfQDIsQT1H34wxxWKuuf8LL
kxI/xKOT88AyO3OSpN4dHIurYKU+bVcN/EkNkhzMbCOfIRLLdEobTSAreyPNQuaqzELukyX2tC6w
+vjnxrUv8Us6tjNjy1bHAnDiHYelcTZaAZ3NRAqzlE17sxWKcM8q//zVg3SKTQ3bNzVAqxBAIOy8
RyV1ggjEMYgjFU/pbLsc3Y+7i731ysL5fIwwX/5Tp4xWExja13OiMBOEiFaWGPJR3ais32/UduyX
ipq7o+yulHbcGvu0W5zfx1G3qKFKsXi0SvzYQe5S0i8ZhX3HgczVJYT9C93pvKLZNgI61B0lnqGQ
Zbkzpx4HoI244sQK16/no+JJ0j23m5GYGvOlIx2FPAgkdrrOvv6RdawHu36NNekt0Jp/M7XYezYe
dCkBddt5BJVVEVjI77FMFR62vGPd1HbjZfxg0b2KZK/BmqESx/wNxGSVunMPY4LUyaoc90J0egzv
wGamVSkujE36eO939jDD7B/Bdn15hNLvPt4lHMy/sg0EE3AhHQ2Dkdti/Ge9gLaTEJ4IWoIkxFKj
gDfCekVeqhitezfD1XbZEAElwS62WOzpCHqR6K8MON2OnE8v+LGULtHlebOwI77Uoh8WezK5uVrL
DGNqPVrU9JBq2tXXAFCEo89mkybpBbUWhXQYYX/3xQ1Ftz0dc6/KZVw6M6qP7h0vdY1mc1HVH71U
wHtLAFf5eVl/g/6h963HbVwhzG8I/4wJbuN7j/MeYwNaNFJE1ps/7WzFXo1c4GxRFepdYjxBhFd0
El4V7HqZM7EtRhZm01FfPUvCWmCl7nNWQd6Q04op0E7NA5Rke0qe9L2K2VEwt1i8693/Cmr67Zsg
iAI5BkcVByrir4DZjGup6SHjm7ZpRzV+iMrvjl+6X0n0jFZ4OgpuzWg9e9Gg/NDzjOX3whp8qHan
kor2HBoetSSC+n/6Xep1vFrpRKA/QLgailTqpzM7nRLwK8csbhkZJs93iSQEymOycgBEXDpp8Zmm
G366CGTS57t21A78SchdecduRQ/9swBlTbV0UuD6wi6RxGUZRN6mc5iPCon/PtCVdE9UGCRYrpc4
BAPZNWOFKGfXrqvZ8nIcKSG1IVVTIbyv+BtoY2yZxZw84PU1I/vDm7igfakuA9JHac8TFwF3JZdR
2mEihrFUTA9SrUJ2AKuFSANCu/yqwVDfBodYKKX9QNbpjsRnUaYYnn6RiN1K4LCktdwOhGI+jnfC
/LYLtqqoGxzG1XCsdt5RGsYNq3X0LkLNBRz4ulZi47SNJKZUUZNHTAJaVk8atObGVRXHmEx0vFUc
jqHgnoO5yixFG8DMMAzMbddP7aE2VsEq9hGxXqqVjXg13tB7TC7Zq8/hiub513xUcEfEmq9FoNvY
Df1Fi2xgcferthT/QKOBJBk3vg//50H8titaT9aUSvTYjP4eZAdEpHkL9J36ztiwDivzkqVIK/Bs
/02pwNye6KTg0CRsnzHxKJmRvaq/bd+gYA1Br+udjrGcZiDlmQPwRZnHYLGFMwsSDHtUk9mwj59i
fCTMTpu043QOFmeEGN2cYO3Ls9VTAhX/qSDzh7MONGxyNP5BZDFvrHspUBhK+gkWbbLrucvAnXys
3cRFtr79SreGAbRDf9U37ibpam2AeXxQ6yk2VLy4386MDrMP/DJQh3JeDI0yNkvOLkRN05Mvigxg
I+SMxRa5jiNXIgxWyKk58cvI7pJs4K+D7ms4L1vkELfQm56jXxOaAarzRA37c96jG+iXIG9jaBbQ
uKpIqMFRE6eQHiFavapa+2eFWZ40yq/mN+SS9iXn+72RU4IXOwbWDBh4xlmTq+HYpXxoBnGK5+Fx
YK8vBdR33DY4+vvTAyQY5kTraPuSumqE2iqqmvKMikv+pP98UlOBkktaNS1m5mWVS3I5kfQHWXuT
eZxrGaR29oSiBdNPrhm2uqD0KI35zv2bcSn3s7AVXhPQozxDrUWwIms7kNS1+X0CsUKeJKaqlcjt
DMmi+XYILqWfw8Ls/NmRz/zxQ/CHv32kaWUTOb3DNaABKn7q/ta6xcAeplbGsRxrD10Km1t38YqT
3i9XtcnlXGVeUO+9iNByKY0/nEKZYwzRJ+VMNOVY1Mv8vq60HjfUx8zxWeIH6W3tOqDAVoMQX0yD
JOrnlD61+oY6oebF32lwppubahXShPg44Gc84FmyXdPdoYm5pkRtIfH01L8lGnncKQxYL8GJ1hhm
fhQe4m1vmoV5mAfHWxjxIcnyU34gREuU6XEiEWArU3uIdb2vBOW/kiGRyTqBKDuqBqlYQEWo0Qrw
3ZKR5Y2zGsPvc7/p/IkPTVJZHoaUncJ+xcaqL63dkrbcTMOEDDpAaa76ImHvmtUnSxC1HBuNsjW3
aA80yviZ56y0Sl5w2DMZn1SWLJA42ILFIJ5bzgX79olPOjBFtwmKqxPntAisdPKblWvJ53khQkHa
NRlZLoUeY3wsNiFi0fB8dHiDztbEc3ApdaoflS+r84H6nvy3XwmURkoaiUITQdot7owrZfG7u42q
GV6M7yIVfIyp5eMozujM8eGeOBo8nX26L51vtv3Jfl0dtayKKLIKlBlsrcWkMVP5CiNQMmpjjxPG
5zD/I6sZJd3p12pbjODT1v+c5sN9FpY/zyuNKUD9HfGvZ27T4PNjtD994NaTL8EAvjDVvcpP2tje
ZKxpGJymoBajfIqq3vzdcW338T7pA5XmZTidctjcSti7wh1oO8XHhMfew0lb6Uf19DYHY0+61L9a
kuTr6suRxNBrmWd7W0NA8Wnk48/ZnOkWzW2ckpdaMFvtc7r4VA86Cvp4UAkjOpQWHQ3hs/vAoKHm
VEsrWWffnUbPQHvI4bqDsoz6SoXBqYHK/YX2YjxGu1+lteiqd6vyv9+0KmSU2EKipQpnEpuNJRdQ
Ls25VS1S82zC5AY1/5bud/Rhiqeg0l4gm6HDQ9MwOpGx33wkrupjGAQIzjxV8Qzm7TqD2Er5hB9s
W0WsXw7uCeiMArU/KQSMCVyb2j6304aRMWe63Cd5T+lgFRuhUiulB9r3jAEhHZGOOzMO15xol44h
by+17X1bcDvBLNWaF0L+GtEjeipevezI44ESNRqMaVOKPSPGNarFfn8RtSNKLf9H72JIvidpNx+x
/H/A8G+zOzB1ciBMYu2cpQOE0b79fvntySZWi2Wmw9X9Wn7pgPZx9ghiRRH9Flnx6FwOeG1kxBhK
EME7bioaJ1lSm+DyNaWryj5b0mQMIiy7T+G5YRF0yp7cMr+qrBR4YvSwe10pxiJUFNjb1moo7izg
TCyj836vRfV71bp9gCJ67UuMfUwFkc7SxmPV3rOj0zlK9eQ3HFcAIuDk2iT1/2oYHzsI6rgzNZ6g
J3pf0UUfBKVuItOD2LZOJMvlyKtd1+xoNMgnJCOr2SGMQn7qiQIwmeg3pJasSV8j7gJRfLwfiEnt
9c7DIfyDXFqVJsrHkYyye/oc7n2sDNUceTq0r5KEcUzrEZHKMzGlNbJHSiTb2MBEm6SL99vzzk8e
vN+cCUy6mj+gzGQJCHblWvt0TB+SncH/tV/Uf5D263fmVp5iJ2iltZMXQJHMQ/DdA1hOD2ODtmCM
lTk4pqsd1AcmefWSm7OI5Be4+oLiki5Kv9IufGESP2magK5DZUepiOLdNFgMJpAgUK92GicqqYhA
nvy/VNTPYH7McfVTdhjsCqijgZ6I6svh6/x7kklu9huHcdZApVVjnKak3VZNsi/0ntoMWCYxLKRL
+SC6D7Ixrgpy5yoLY1QlExD7/cfOQKBuVyTIy/C1hXmMrDq4I2a9ln/sLzCaN5ME4wsXv1lPJ+Ij
tofHjgr3QAsrCFxTv4gSQfenZh1KewvlxXAL9kznhD6ARuf5Xjzk7ehTtlovt9qWa5i/mb+2I/mv
D1ci0Va49PqEfon5y1cLzDNqLwihyapbpvVsccI0GyG9J7ltX5r0DTt9kn9cheab6nwunFnAt8Yh
ogBPJH0nLlV5pJBoCGOfIf5Vncez3X9Xkm01+R+1R32bmR8vgLa5tQMLwx5cvVUPb1eDqNnVzT0R
dm4zLeV6aB7T99nqjr/RB5X5LA9KutwcUjQYGV2HxIKoFC5e3/S6N6CKe0qLAco4yj6qNKQa0wND
7G2OPUjNQS9P/HCQNf0TaZ646+sPigdwWMXR61mU3NXmmEuV/ZduM3x8Eev509tFmCo7XU1ac9JE
42kQpqUtIAaMM8/AVkkNph9qgUzvvl/GSCyKumPxCztMVzHT+2nHEYHP78fZKjfvy8iO/EU4Dqy2
2rFSROmXanY1NjRVUCcFMSydJmjMXVudQ9MDhfT9L1DkaN41aop3Ye2NmfYsPvBxGiJM/QFZJrKW
ePVfIiWvfMiKoiixQ78h4pzRYTv6CTq+2t5usWLseHWCunZg/RRJehldTWkxVyeFSCdm77WhKfYR
+D3t5UhZQO2ScT8rUykLD818xxSNzUKxZENEpuQ2zUJXjgbnKUxu0UqiE98DMWX4N8lHIfhftCIY
6ZI+FPIQpjdUkaVDHl/cWwAatr+v691+dMDmFmC2eGtbtiJOj4UM3VF3ACq70F40jivukO61bDXV
q6TbxzjTesG897ZuxKrVqgC3OshwXzIgGSg7bYNZExJFLp4Fq9EgTyt27wbO5ug5R1q7g0qYz7+e
dbfFq1W4SJE6JKpRgqXn1QuzQdXBYUbfuVzoCC6QFNRadQyU3NZF5Za5PWTkxc93p47jaRVtU3e3
c7BOyu2BHSuX/SVrjpfzNH/04b8dUIDpUvu0ptJGn2OpQl9izBUoTea5hJ0qBZKZXS9c3SRaYNsf
rZEJXne54GVPA1itMSWBRDyUYj39BogkZgzheMHhkVHh9etOHN006EM+NKmukMsJC9VkIL3/GlRp
JyZT2qRl/EX5LyfR9dOllqoquOk7/lD9sGmE++2zN+3zH3eKkj5y/FCKRySvwXDQb+uPx9oAnB+W
3Fg49vK4R1q/PA6/LlObEv8u1mb85vkak0/2wm+93M29N0Wm60pgdQFf8JjjPIVkh/R+D2vLAJA6
afQP73z7cpDjyxcjq6QLh5dSFH28O9fg/jAmNce06o3/oUChLwYbXaFPH1pY7V0qyhfFLvishELZ
HBEGNY0m2pa69rz5V9mCAQJFUbGum0hw1Gh+e2qyVDMuKYIaswCz3+012bJrQ0ug1Jk/RZSxVYS4
o4f78a40cMx/Qxh7P8GPrpl9zwmUPoNmRzcOlDRQ92YN+4oXx8fcVeLXnXXl3hVF0kO8x2BYoU3u
DXci7IAXRg7fmkutNO8QziDJNYYscsBlCUmqnqSLmJkd18ZEeJ1Uze7xD8gYd2Ck1HO0ATPyyK+O
9XdByfsR0WOTOVArsJvbi9ZNLb3LDVaw3IpB81IATmCUwcKeZVO+Byp9fQg9mRZckm5bRsvpPCxk
Tt/lm1L1t+/CsdlmCyZLgv9T9XCS1ZxOIgnvgE8OL5YmHxYqOwbqqTlq7kwIXXEOyTDpqOqPzx5r
RbjSxp1L99MLXhkSyN0/ihPTU/hjibxXNx8eEH67HBTL5CnhtN3K2en9dojtpup47a6DOB9KoOPq
+OkTpGZsidkjguY0GB4qq9VfTDRVcUND3MtThMPzS9Yv/u2svtcQVw5t81femD/435ZWu6NFJKBF
baW3GjixDP2HMorOVoUiulvO8xGSQwzfkcZ/aTTWqdsmPiQwTi4Lqwd2o7aKeG6/WDi7xA2jXmNZ
FM0t6h18IHY1zsbxdhGueNH1M3P+Qj53RvIREYn126ACzf7rbCwQsnwKiDhYB42WeDYs0VFvmxpB
Ua8srQtL949ACnJ4i61K/LJ2xRAMjqcyRys+8sNojhsA2VKhyuOzljlqoukjpB4v05O9RfurfT0d
XW8g5RnShbABX5Xn3vNN9ILjumzAnyspLmY6sGkkGDmY+4VwVNwLQG6SeDLOdk43iv8aPJYDe5qk
3g3M2Tbf6ubCffe2J0XWJ9Jgw0JTHhaqRAsooySIfSnOj0E9VN/gPRTqMAXx0lcaMATNJFMAkV8V
ueq9O7MwqebzH+aswNMtlDY5f+TDjYPaiCoK9Z6O57yD2JZFTeECSVgm7ERfPEP1ZEnCUoboeMiO
2XdZ+lVLEd3OL5VOK/zSvyJnM5qRWFozPYuNriIxnAsMj9rPP8scmJC5OESak0Mmb9hKE4J63uFH
rsN3QPGnwArsZV8tXxog58nkNsoslFGAhoDESXW+/PQvnD/UV/G4JsV1ff2xrzQtbBljlyrh+F3E
qB1Ijr8zSyUnvjLN3sDCGDwXlxjHDS5qEXRp1Mlt2ohjQiud3lwKx2z3oNXnte5xAHQTXeKwiKxF
RB7bo66RcSOB9lRrc5eFvxrMnrT2ENtxB+b2z26fQmgB/7zM+dsR2vpoMLP6GhgQjyw37VgvOAO0
Ass+VbAyNC0xXfVbFajp9GrswSOLOpoZ+x2L4sBATP6K7YbQGDeiWGn1MRIxz/b0GTXVE+poelUj
Y/MaXKxDLOoSpFD9UtnaWcv44/+NY81z6Syu4HTGeTm+THAENwNaMZCL5KMb53Fb9wgZfJthpnRs
X960Xb+pA/ETv5d9r7D10NdfLl448Lxxs5qk9NWmZ6k1uao8/Z/uq1s5t45A1m75fsrwnMOiFKfd
kQtiOLc/7SbJcAS3k1CbeDgp0eb7f0A8YvFdFsN4qvXxiEQG6Br7QpyBY9i7n+meHFQrEkhfjOBC
sSCcY6RnN5SqWnyontG/9qAQvZXgc7sjlbD4g4U3DBH/ly3XY/CxaGlnqvHloBRL1qtC4tK854rw
zsVwOcGChbDchFkjbxIRreCSBN1DTPBG0tltWE+r6RA2nq+qMxXFJvA+i0RyU7D+o9XR8mX5F8fa
unvH4tzOG7E1nas94ydwTRwMaRHPHz+iqMthyJJf75RKH95heIETPM8K8GtnMZQF8nI4TRBV+rEu
Uq+wDDBvYffJLFr2HoipYxTgun5WsiCHfxEnIDXlfse3ADwswL9u6xwLTM9wtnCUyNBcqiUsHEfl
bEdmYQiE0jMl5Awj/2dI9spXrpmH6VpOVqMHS1Gw7GDl+3JjHZhGlTrhWNelpRvgKve3uWahRhgX
J7dIWsZ9g4+EuZ176EkFCAY5HRyaJb0POStgiMOM0LVBbHuO+LAsXr/HZGLrZ57MoQoPzXVk1ZKG
d4VRZtj/wB3ZDxUzYXF0TwPaEJ2qmDIE0eLHavg+cmLe6ycVUkS2KBkewzqyiX3EkfJHu/q6C4RL
0lBtsHOb7s8rrN3jWp35Ne06cLOdPnPoqgAf6r/hO4DXVobnDJwuXW9WUE/e6cK+FsnWnH0po22y
brRuWJ3tQEeSslEN9pKDfJUmZzaL+z/yztnji0IL091qEPQxfLFCLpVJCP/FZw3I8qX2wo3yW6Dr
DKLmLhFyL7HZXcVIHkUjsXMshfKEosPRb1C+X4sv5LLBgQpihYSHww7pYn9uKNOVyclI0i5tDXiN
lu6wQlvimFK0HP3VZPIk4fhFVeEg6b0DYgu7hAqMcyZd4MSEHhtrt/hkB5bgoT9UTd0iqAmgpRW7
NoGD0xCuVWeua71pPbjNIITDFXi60PNwN+9LF7/+8dkH6I5hv79vo0FD2bd0VdNbv9h2fjpj30yM
DJTSx8zCqoSYhk1a2cA7SKzU3T0QzUfwIqgf+l5s1R0L3GctzUCt2XFgOuUAcZz+RA3Uud+4SmDZ
HPELfel/EGr1IMWO+k3ub1QouK+xkx4uT6QEkzCHx00jtmJVTXTuBibvcrjBop8lFGMUF1mPrV9H
3Al+qaHPxDRFRA3xm7L9JD4X6sr7iFJp9EoMdJSKDzLDMxKM7SwvFbnnqFb5rR3r2Lmy9k68uKva
VWv/2QkwaClzUC84hYtuaYvuCBWdJpca/U+R3jEcgzvlDNA5oxZRAFXsHw9DWq1wVP2hRFTabNoW
MB9Eau+STUgAfbuVQPEbl05YJlanq2K/UGlbe/uuaonnIp/UOn7u6Xv11+dzAUBQBA6Vt9222YqB
m4qO2WsgGpRM/sO9sw1drf2vq5eP0/xILPhfVyKOEF+YZ3fHW9BNaHiAZETqm5RsHNlsy6OlDW6I
jJoNcDTfzWWeHeoZLmerRwc2VzliKMScQ23ZtLt3LIAobjQvVlXfA71cOHrlM6lcoqgnTXN+24xk
PRAa1xIqJ4pAoN2JY/MWceahP9XnyoeIrzJOcrzOgyPdnPYv0Tl61MShVex2zlbij6A1iiY1zchO
y8nhWmBwxae0/CFZZsLBJ05KHVdFzMvlUYlGToSS+Vs1pJYm87cBar9U5EyPMxXi0XjQUnH1kkyt
iyFq01/Lgr1bPb57q85S4ZARwCvH6o43/wQZBg1RI73vuhPSUDjv66UlrRjD+pYAv6A7rq7pmUQs
S2vt2PzkiVwfbAKSRn47aJ/S9GlbN0ktEeCAFV/PJN8UDlDGv6P1uEOLwCs3E6lthNbajVTjcBtN
KF+A1uNYaheajQK3F5bP+/4jLcaWIYak/7SHjtMXIE8iMPVcwoKzDAPwJlfKud6xzkfBBwcH9PPh
A+jR0Ysd1tOAO7fmhFQhw83pscGeBuqcgH76UF90TB1a6xV1rTsPFsur6bOZnzT8G1X+T5FePxqp
j2mcGLg27QOOEDKFTj2jYcRz7fg8KppJ9zTWCDsnU2PLfCPV0iVS8aLyjKXtTzMa40n0UuaCzlAv
tI8Musyqtvrgtv1/loExL40FET9s06BSs9BNWiy+g5xuz3peaQVBw98xijSNew9iTfNx6g4Qqkgw
DTwrzweJxVmKjirCffd+oSNmC3vlwn5QYkDiblFQ+cKkEjFIYFhuBCC4QLKVS3ne96m6fDfFSUXo
vfdsKynOrurL7gLqRtKC3Y+4fyrLmpYAPa7+CT8baHzKZOeZEcFZBP2AoCcN9aHJATJeftloPH8e
2Cs7vrBqWkacLBn3dW1MPerMuy0lXa1FLj7gsAJ26yCZK2z1eLigLkIQqhs0qLPcyodLDT9/3dbL
iQZi/NXcYt4BHymEF1iLodkcMUQh9JO4Kfkp3X+6QxeLLwx+mVnETYRWfnIrMjxoKJB+/CM2eFQB
K2VPH7pQY5/LKnVNzNlX9HVV47FYqX6qu8V81TcluhBhkYN+mvOnrJTP/Ka8fOz6xhf0kFit37wy
M2iFaVgqBkrJCPJs05y2iX/uHhu9FuYafMItnFL9zO0vcQZPcslFcH6ZND0TrJbSpSJjHPCLP8pF
1fCgtPRlH/Rmn89f7Hl2wjYJEdW3hBwy/JLB53QRspF+AteeG8OT2k+IzQHAfArwpLe5Cs1kL6mM
BryOzFygKi9Q7QTiaIisr7auVGkfEZhg2cKgJUnkmcti4Dtd2W4IE5zfGB+OLO9/hE14m6hVwzz5
lsmdKsw9+X70FH3jUlSVw/MgbjLPBv2TXspzDOwsluq8WikydQUwaEO9G56FI9Yi/hqZ6uphTbCD
eLInuULjCspGBlMd+SXPe5p+4gpO2RRe5AJtI0ON/1XAOGhFLeckiiHlL1fHJvmR78Iw0thdNA9+
IrsFXPUkydMRFbD5LMP364+7S3iV6aL6cYHYSiDm3odW7vle40n7jbSWdypOjLhcqgeV0ARP998u
3MUCm30Ao9ZphI8E+MWvGXk4htlVLEk7MOGEz9M8RHlqwVK8YNgIf4OZSGWttH4dKne+KtgnppjK
y3CYyVzPAD4H+Tek3K4sP5N4ndenMpIdp6toKEyb+KxefeY1q8aYWniI7HmbkPykSUba7CIYDrvO
RLYrOnq3uXxRspbTv6WZPjhXh/eO8F9JeuP90jPhITo6LLwdNqG/Zfg3rhicAv0TVNZf/nDGTmq6
fswTRswOcajHFa4aZzlQ90XFsn/m7SaOOnV6dJR8Cm963nDxdkq5p/4aHzs4tVJ2jjYXHcJm/eAz
XfwiRSkD5g/Y3UxTuVpy838pYl1FKWZ1ErbDARCyyzBYW1IUF/IbrpxiEtdqvYmf5c8z3Vs5C8tY
kdtXiGWZS9CC/UE7WFs+6s9P6zBZVJAEk8+KEBZTHy+ApfnYSkjwgZmxx3Ctc0XRh1OS3qj3P5YF
nzS7+9OTjRQYHa8oPA+pgdXS8m9sLysJI13md1P7ATsEVaCmB5DbiOGhEYha1URjVbIqiwUwnZWn
QiGvsqi+Gv0xwIIyt4KsPIOcEi1r+HHXMJwgU65mm2/pWZRCpYpLGeiDPxQ8mZcZkgpAyGHTrHo5
fHEn76leDhx5HN07og+wDB9Z8FSiuaEW1TgLXqVbdKM/s8TPo46wAS62FsVM48Hg1lW2bTF23rJZ
2xPlbvaIfwtIAFtx184VweGucfCvKkc7uMfcThVkIorz+scA0i0yIegMkCUYw781QaUgiKYuwV23
uqnTscN4+pqNdpS2RKaPkEF9MVotd0eWP9gxbjXWzEcWoo8TkvZAhtYQ0Flq+pvU+IB9o89oiemg
xC1XbvtfVPNWa4/ynInMSQKOZ3v8SerJYLUStvFwoo405mWLw4cHV6Jhjt7HrhdvmVaZ3gY+kLeg
g3njdvWhRpcKyOA8GAaAXBvzfTkco4FVXRIUcv+0oSoRwwPmZlIgFDmv05nllmvrEqt0v9y13Qaf
esAKiahaiU2ghfiItWH03gqqLhvH15/6rLUAaqayGjWb7ABUX8rQzXQ0ZZeVxghUCmKeU1y4tDj1
ONRGGyDUmmjQZWYkZAnursQtDaRjRRYndS+i2fRaReojIaHVN50PhL6+l6UMMGU6TaVzPUpnusAI
rxvejgeM7skMHJR919txNc3rWNhUMm9Xtq+QManNtTj634dAJnT/KBYdKsa3iGehswBWvWsGf4HT
QtWbh8OOM3mGSE8MrKA5Ay60UVaZynnqXXLHK7rNJL5eIclQ7OzSWbxfFy/bIF695qgJvIkt5s3e
8ijQHMAK9DlKuHCdsjxFyA0yChS3DLAvQcxvIX2lRowgufRb1Com7lgrierCozhFTBHuCTMRFcOa
/4V+NNSLbs7n3q8XoNwH5yx6kv3evnM1ttyJzKDKGQPWmEP5xBsFzCiOfnomw2kyaTiLTXj/AgH9
yXXnV1uEMPK8qt7KQHAC0w9Q1zUwG57W9RznWo3fHoqR9M3FOJcf0kfcsfv2ASyQUnWVuzkom+fK
0D65rHlgglOdxLQAXrQ5lGLVUUt2VihUTfmKmSELXOlLrz2eRjaiRZJ/DDT72BXnJwShAhI4UocH
8DxOQeb+SfKuhuJDHk6IxOxzp/rvtG9fKuX3S6Bns7pq+8unTsWkGVpk6EMR2PohpxaHZL0nuINv
vIhIUrG2UnHkumqhk1jzr/lo+ZJJYJqYlzmxIf/QJcT4UjnSfzwREh0qSbCG8hsXkRTy9i1o4miD
EJ1dgnbVGIxGSlc4Aq6gXwzOHwJp9ap1mGQkl3sXh+HIvR937Qf2BNDet/6FDXOpzEE1NihnDuwy
FXnZjZpGLnzJynWClduOgmJIDn0xr2lXlH2Beh3eD6LwORFZ/JhdVMzhtiRxNMsnspa4ih77+U67
AigFcVaJ6ud/fjibp4EyYlYthq0E/P/RJTe2IW8t+BapyZ2aIvECWrPD0lg0uszYr7zU4pRxCDmA
DnXRzpM6dKECZgiwMbaEdF1rWKXYN2bECSeRZcWba78+TWKaZKXRA9a74BAi8qymT8xbZVLVF7iA
om8bBLlUTMh+GYOjLXoEkoUOpEapNYxKkLvZyl1qmm3V4owJ4fxP6PMniZpbx+QQGtMgxN4+YQce
0KzqEDV570NH6/6Vg5UBO1OtVNqwH+RmdMx51mkIS9Ki+b/6wNw6j3IGShpmBC4t96YaGrPpOzZu
hRNqLNAXXGpZlO9eXMb8dASniPbTktK+jbRPtTvXH3+zOwRsOu6dIiuPc77sxiw0bEeBcuKIv43M
FBENTYcoO/CUf2cITaz4oRGZjbPcn7xWLtcOiwfrhbRitB88yTgOYMw9NHaHAjxtiEEogUeluAII
klXwKT9Mk1FCZCtQuGvTu9czFdJVwagKZukgDwO7yrRF9J+5AyK4wEr3y3SWOsxt4UTBo/MSnepP
BA56lPZx4jtfsdUDi2glItAAquzjeY0o69jn6pGO81xJdMrj+BtnE7bY05bmsfFirz512W7DEba5
gAE7R1D3qGBftrLtRuRXHAPCMwjL48mAfousnwPurugpTeJ4Rou3LtgE4CP5ltlKB3TQ433OoQ1w
vkhmN7Mc84zHmzGhQyv6N5IcfhT5CwWRDzkCZOEYt9sWzDxV55SthN4cPtvORopKnlvzZv5tDE+C
ERZZkeyAo39fnbN7OZJIJn4gTpBrN4kWZQQ8MYVklLLfILy4R/g8EkQ+yoC6Mv8LaboCVJiJbW4H
koU34Uh1SVmjNnkH8/ZQQdYsqqETh85/IqhrqE7a3WGDrIZ45NKBZRaG98rjGBOZnLEWQCV4HWuh
HBkDyzNfznURp1q18F4QOzMncKK9NVCchccedxpwqyU1xmYnPhoqbT0P379w2y4elFcEbGZz3LyD
Xo7KPxPtO8PU1oLUTPxKhowNWKpEQlafVFyLxyEuKIeKEf985kXLyNxWrGoqJE8J2TRbpSxkdY87
Ix1Mmc3sRNsBIrg6Yd7yyIf+8lFsn0J5JhglPYuRkn2xHcCc6CfEu3jsaKhVZKP2ydBYjAM7VGF+
hUkXxgY5UhGq3Qgh34hVzcBEaiuRup+wm43yqho867ylKlG9pSeKCrKU02GVsJHBy4M9etZ0XCxv
x8S7+vydy01vFGqJQBLyH9DMA2vDb04zO05mLjftXJKoB49+6gNg3ua3X6cBJA6vEJubQtvNH7lW
kGVdlFLEV2TNCW6SYa3i5kDvgXTLaIFHbzw04g2Xg96Vmxgus+fyu2J6sMVUEYnhbK1NRWlemrim
Plec0wV1f1ykBpWeJYgqePeIgkOhEYtqsWgu8yhpiXI/lzGWd5PDwmP3K3o16a/IkEOtlXx3bNE7
17uGc7NnEb5Mbkb1CBrZrCV3QZluW3/ivWRW8GZkeK6ekF9cZRHV/0OtzwZWeAdrvvlInj1sCdJV
BuT//+Sp4KWkh0UsrYANKmgHag7flhtY7rt+2LLoQKQlo6ZAWi1BhTaA4jskOpqwCdZzggP/33Pz
6bfMOthMGcJd52zAuR5kf0+PNh5A9XCLcUQvAPLhzKzihTEPMNH2QIZ+CzHqMYVJF/clK1pXeYHr
7kQkhlZVb0HBiXjS7v1lKdr4YobEAzw/gQK49YfjhH6CXuFVQWNY1jYHbmGOyMVZvDJCl2bqYAfX
XUcgPwb8br9uHM6kfF3JcEE2mK2FjUwCWMCuaAbc+09RukwHZIOcJ+ic6nhV2qUqLaukmHfUhjzM
2cpImJSr4LagFcbyEZHIdolBieueItEFvKnbETGxauAzDvD2/oJvHG8DNchjoLSceCVY0lsrP+Wo
NHKgrqhGirC4tikA8fkx4ic+444At6TNM2YMuRXKi00KZzpoHithtucH2futfyDYEUx+hmjJUrFU
E/N5cJMtjkFRKMb/zefxsk4f8NknxWCHTRfJ/DA7UveNiPRpfMX6AMEGcjPDbV5pvKpzZNCY8yZj
hY0pyTEzet4vN40e3Z0hNIxpc0seYocaI1ktkCgtoEzP/GoDHpAzMX8ZRNhNLMFOJk5ub/mCFazA
6RHXuqUpb8lLQLs+7637niPbBpZdqIi8ojOuxBiw765cAx40xZzJfefJcRYo2Zl57R0k+ECCJso7
hr1JXmgHsS0M29xtH3hTwXX/aPs3RUCEFlB6shblFuMbjwjMqoreEjLEE3HUgbqJw1pM5WXAK/Ao
4wdEcJxu7MMWtouMOMFEuHzX6eXzUCcng9qoikQP/nXVNgxN9hYf430kT52E+JzTh5+Ap7MYr6EQ
wLdtEiaxzwbUS+0g1Rvat0Xvy4Spt9AY7Si3tUZCncbDQkPrTbjWtF7c0IXRn+F6MOV/9T1yTti0
eD/3u3QTju1w/Q3/dWbf/YPgeAsz3GoSJmi7XX07JKdce3d9Nlt3FF9ircLcqKQAzn066xZIgvlG
4HVemQIvjF9RELY4qNo4KvsKWbElbTV8Kj/GmxRe+SXTXnJVs7MiViCc5kGKqHrO60URF/QhVTPG
SGQuV8pmgU7r2CEFIayuGolILv38c4SFdV+hxMzhyy5ik+M8wzAZ/7F0XDUR8CUDL8Kcbticpb/v
MFzv6BpPEQewpDNj7vyRBbfwvjq7yhnEv5Y3eRHEqxuyuEpCePiYDiHV/1ZinmxxitjXUFW0vxVH
EjBKSNBxf3gJWxdeG5AJcWjwZVrd7oLXjPoPNueBAfty2pkNwopi/fMcJuaqx4gCtd522y5i+7tO
/uyLV8mtSYDgvW2BBC8r6UYRNL8HzsCUrtt44vrzKpf041vuQxICVxmBv1NsvENn8MOCckeqlTSA
qc+AuARFoR5QLEWHm8mNU9rTUkcpc5gLOvX6BvGDxomojB2VeGriAi3rebjuYPHfK8KRue9Oi8u9
U5FE6Tx1NweOljJsHk6EzrqNhqvEvflmQRU5rYMeEi9QpM+anIcJGtWRfeuytienG6EDHzpmWYXc
uthSjep6a2gA9p9GSO/ihBhNOWQReRwj87BaONrMg45EkmJga6SkztoMw48qIdQSZW0JnR3o34+N
sOIirgROJHzI7E6lzh5/72jPSEpyx+12XtCbgvrexg/z873HDRU3cdoImR9dV761XRuyWvUtf4EH
zKh6AiMi16DUKmKQSzLILaiih0oyWRC105BiudIHtAj79mZEgKM+3+oUFSV+N373XvkCAdmUkZt6
ZYrciM4ANOAW9HuPtJU701ljHWOdcNE92/pCNRmnkpBiYnSWfRCYEWJa0/888yRjbyBlo/D77H15
7DHz7tz4vzNqDOmkSGEJQAmp6zn6iIKgCGRoNiYEonGIEFaN5N5kqQdWWmO/CO3+Hk0hCrxjW+Xt
4aXtRgnIOLxD2HcKS0Jtk7gDiZXu7/zUGBYsvhjWRDMeV3SjEy7soYt1xsTGNUNZvhFreBNs6CO8
eeVoR5bQT+auLNrufCEBbou8umDpXuLTOMkz0frHL19maSlBYoL3nZBHZVhnMrdQgsi+Xz7WmeWK
M7ceHMW8xv5bxb6BXBYqcHwpeBZy0CRSOjcwmaGOCeJPOV9P1scyeegcl3up3t6LSKFr3xnu7JPS
Z+NyHuO3C+zTIM0ZR86p8OrAP7umma4H5kKcs5Xrj40anOIVDR7QFXfVAJ6DfZpbJb60Nditvh7F
MQuFN0J+yc8L6Ned6xH0gY9vILE+le3HFz56K7Vgr1Y0XT/fDYJi9qkhGcIuM1hnXc9dROR1r2zx
m9S24KCwxGrhbrSynwv89OuAnck1o3tlstrq+6GjGsttqY4EkFkewl8tEQv5bNcjSP2GYoL9ZAwx
ecReiiUewnWgqUHZzda4J+s8AZn5Sezo3aMR6MXf3FgUBcqJPMjQuP2KiqDKA5jZ0S4aelUL3TtX
daaucU7izLalOXld2iuZnNcX4v1I1p5/b3OBUFLKgqxuwGeQ4dmLwFyWiEQ5p7F4rDSivi0Td4cC
AS23n4mQOYgeofWYotVhoJqI1ld74PU6PxrCmiZs6KAWeebtCw4qhFyI2eitM5cmfiWKbH4oEaVY
j1onMoWFmyqSifWpiwH6K3Jek0Q5X614JFyzYx3mivgWZl2gnt0zZfCV+uzuMJ95DrdOJBZmMxqF
g8yuFFaELzP90RHEHMRPCbpVQxslzs9Zexv7Uj44p2vzyoqfFMtxvyEYBTg92zc4jyLN/5u6T5Nq
eQtlbTq8aQPhOUJltBkevZ944e+hIJtkOGxgaXwGRDqS9lyQDMPv3yfOxdvu3k/Aus7EfXRB0TVT
39HVr1S69ARapmc9mZsQOdPYbdGrtsgDFU28VDlQDUvVpaN6h6PhU6p904rqnjtH3JPLkYMiMpoH
y7pKzeyYix0vIEBWwYKONbvpmEL04ugeMpb/wR/32zA4AhVDq1BtxIgIgsTwRbE86mXh0bWB/+mD
yeyds/cum4N4quuln1aAvLLBapZr5fpdardD2umiPDZwgfRTME5Xb4/v9+BKMCiX68/2FyP+ocv7
1MxfIGeUtzAyl2ys3ZeXf3/oW7XgRSli0BnBt5xj8OtFME5qOjOOSJDCvRBTVcJs5u27tcYyXOPs
x7ZlJ8SQ1MtSRg04gpvglClt0+/zPBUY8ez6JRK9YbrKw4/KbMf1qSX33/zD+AIeIjla66rU0GMy
Z1mK0nv/rDFnRolqRm869h++bvWml5K+pOVbaZDOqKsuUoOlsC9SWoIv05x3FWl0GkoMXmiPE7Vd
6kGRAVhHuom0ru2k1vO9DpkGa0ACRvi69quuZCXzaH1lR1lURkrEaQ1h9W5RLxPdU5mTFrFCWrQ2
eXZTBNWPqXtOpAIMOuPmqKtYJvSI693q8UCb0yyk+0J7KxRglUw357Ngt1DVCf09fjKxDKHNmoxf
n4Lj95xZbKBu1EBV+2zH4NSfH8ynIERHMNkCN2o/he1awNZAr599bVFHccyYHe+X3sXu3q/GWtAk
nnGp5+wWb29t7aeWPpFnkgGgTCp0t779n+W2UQ+2k7vasXDWot5Tuv//QfBwOQCZhH3BjdTKIca5
jAe2muLoPlIDQN5OKNu0+33efObhN7sEBTs2V/N++IagDXiKCOyhr/w6u07E1GnrepX97y1FjZfC
DJGnqkCyaQ2FebYs/6k3zXZLam4Z/dLG0JzjHnuZHHqNWK8zCxXFfD0dF1u3Q9hJePJuJV18HdMQ
wiV+LNPpGYFbQKEn9XnhpE2/BILoPadwF4OMtRlzqET90uOi71huLTMj3h/jCFof2ozDAscj8XX0
UwfVgMVSlKxObsqmKnkOOIJuQdBFi2n9ThsYhMxz0940T/Npvl5IiArwc/MtVE+4Jk5iPnb71uLw
j5zDjzEvGn1wPsg8mpY3wFxV9bqAO9CxmxLPEoT/aM47ISM2VJhmEi9/a4Bhi5aPN5E+4U8EMyE1
j777iAg8Pz+SN57GZ9yS8oAUb0yl1VK7l6FJ4x603BuB/ObPHZcuGsJb6Punqlx3jAY35LHI0z6P
+pk7iyk8yS0vl//bnSLqX3X1Fx8yQ1+oyTvXQRvwMGcVO0liTPwIoXV7AVHQNU8A5cD/ybQctW7k
2BL8S59KeG0iYw//UqpQ9yAkhKdAn2iNEeofw5dyVJ8HdqJgEtrFJzCrwZRnx4isUf6czPV8g2aP
XsNLaved3uGVYxgR0JKUjlopwS7RblrOSypsDgUDzcejdNtsJKKGkKSO9OuWiLlFUeG7mi9ZdLgL
iTp1GJC3gVSCVMTurBvuUj9sYrKkXRcIOvYHRoXJgM5+PBuAtc5DyCrd8xStHUyLyVrifSz1I7vT
yKHtyJ5AJpk2rhWF2TZTh3TorfL/ScUrZn4d/IfBZJkFU0Vu18sQnKQuB6UbrpYAr+gXEzJqaueY
jZk2mMNTbF0b9rYnuN12zsUrroZ0CDIl7OD3nrzWtRn7D+A3/AAHL+YquKpJRjIZxFvWvhcgNHOP
lf9yIzGVbNwiv/OVAuZQiDf/WrFc/XWEWIYDs/MwCsYAAT6cvS7nTRFo1rYk5ZBHOOOCA958aUlL
fxJJImzy7vWgYA2RAKcc6ABeTOxzQvYciwMQVZHFforNMbMVD4UMmy+TsflCXX77253vYnnlPXYg
0Fg3BMYJLDUIYuzvJiXhPzZKMgk2uYeRXbjXb1KjY2Xg2il0xxsjeorE6vq3i3BlbFgTtBEZuejb
1HHxmPGpBiJ7qjc6hbAt3h4wX9lRja1S/Qn9SvKjT2PSSVz3yo2tv0SkkNzrPF/q89jVdEdoGPsI
8TnCn9i/EPDDec0ue229J7naNLqRrvc3oCMDVe2TvVHyS25dgL9wuZBqn7mikr9zTBFYfWmPpLOt
NkVyh0+JcQdk6hZRr0tkLl2CNayBXR0zqvNANhKX37VH18bNlC4WlJbmhBseASWwy024vgu+oruN
pVvcu99xVkjfWDgdXFCVI1s/vNQdsr7TW0nDqxGrrr4L7ge6ivg/oXT3ppg1hlLFi6NhyP3jJeAd
ueG92M+wwPrBKC46t9nyC8J4ioyag7H3fhYeTrqCkTX73VQpTrujAJcyqUzGLKPFQcD2gaFa9G4f
/veo5BC87Ze9QSgMlrwHxhIQw4PM5ASbCmVuvi7jXwuv5smmyf1QVDhOkq+p8y1cPd5yg1n85Amy
Y39c1orzN7jGDmvXyxWd7yRAbGHY+tXXpQcRiVe2AFGCaiL9rbFw+jtobJ8xOgDTZnua/0xBaYOZ
JcsbNiNPILK3v3ibuCTMN+0unE8cZhfmXzzBgaSHrEd/DwR9WBvxW/zeY791jxdeyc+MkARVY6oQ
SvO2WW9qqA02VNYkMguLPDD+bEzCOZogVd88Gs1740gebMFUPxQnL0o9S+k9yfHDD9tm5rG/uhuo
RInLNvQkMwqhCqqgtdzCE/4mgyQt1r1+InC7dpha7rGs8Xh+3X1h/7z7lVwqX01iGrHqa45t31Gk
wnk0uqTInbmwO8P7yA8YcPulm0Cl4IWVA8drTrGx3xfyXhKRxbE2qBjv8cIX6Zgx7AF1zfBawFCi
FTHf8CZYZLtbFnT9wSs5xhYAZRfF2QH843W8/ib/miJwLVLAaSOS11f7e3OPgn0bah632osnuk2T
BdnBPHXv5nnmF8iQJEUscvuv7pkmXggsAU6skYteOb5/am9pwuvrXlYIzET4D8zjtOXP3m6hiQtj
6NBUpHqQQAcD5X5q9op6RLPizvSaVaPZ5Myb1OYboz+Slf/94lGKBFzqDamN/2HNeFO/Q7gHlZmj
h8MnkzObWczP4M/OdHdfgi0jSmkgvCTKTlnEXEvwQFBdcDojZJcpugyhjPbZK7aUIBvbnj/JzLNU
L8qCpPr3DgKJvwTOSXZJI6wUOcbmnUPZSIrlCwI+Oxaox9THTX/QGWeGj3FkS3I34WHPzM5mLd5j
/c56QkVKe1TJdh+8Luy40GNX+1qAhVGY/f5+DdLRn48ciUQzX337fKraTh0HoasmS8UWVdeLH/d0
PRZm21I04eAiXFBiMEqii27r8ySBj5cGPXO1dUY4qVbaqLPfagv83T6Mqlu/2g+9zQ2m2KL8HFWO
9UbTey9LCg+WLfCWNfBrc2kvzjUPJWhu/o8FxQTnQqMO/4vt9egF8P/q0lpn4jT3vmLbB8NHzU6q
Tl9hL0HWX+GPMmNk/6k9ZAyDh2ZgPPHSneF+hPDzc6TDEe6OrTFeb/e9Fne4pNaUtQuStB4JXXNM
XtDOkcMXkzEwdpqf0+qPYicOwFT1fXPMGQIuza4LKEyohFQtE1D1+BlnRRbzBIKoq4JLYb7XxFG4
c7CBomnilsNJXGIMOZa9G3q+7P0mb0muUK65e5CL6AhPFPhn6HRm/uex5NEE4u6FtPuZtUDQitzT
XJu36p9Uu/rr3v8QowsInz14Ghkfly47FaFmDFkkJgxlCl1j2BEpFEQIDs/z9sjycpOD2TtWapEJ
nshldlu0/WJ06sKD0g7jg8+ylX3ZFLu1asp9GAhB1L1Onbu3AUbeUN0XuhhWIFFjfj31+9t90Brf
HGieznBH+i7u0XNc3WJG83WP0QYi97VzwDvGpmBvtpPafj+F++b7tErY6sWo7CXAu1mp6hlclh09
jgF+NJe6n/hc5ythYb6o93q2KKWTOtLu5J11Y8bkM+liop06IisoHYDX+HMprojm4zzSFMRS0ut6
s5w0l7UNO54ofwfakNYTgj/6ZoMnGatfKhgRlBIkqnHn8LZcboNcsA5X/wT78hTgnaGGzUJm9r8l
WVcNzOqQ4O4wLdBxdkTKvYVnqDkqyA8ySkjbCcpkw+VpDPSa4annFEWqSadoyjZlIfbtoxfKvJB4
BBEGfyXM34pDK1BY6WbkEdpBWNc8g8iqx7IGDp0Igia3IH93Hq2/Q1vB2Y7y5cHmhyLhD+JmK3Gn
/3u09vNBswUt16Zsi4ZkNzuiQEUKzBgEapJKHEWCncuv3WOsuYPgKIDJ/xMRdy6U3bKgsOXMg0LY
pFgOeB17Rwy9MiwSorAW1qzEhwYCEaqBtuxfXWoSFYY75agSP2ZSZqLmradk5K2117XVQM3S59dV
anHb3uNSiVK0Iiq7Zk3ufzLG5BRfDD3+DUHBdsVEUIqCbNWsdBqbpeJ/0+3hZHN4ykqZo9erWPXi
hveUaMl9pOFqaHtM2/sS/mlNN2yLtijqYWmwoeq+rsNIKtPoVlEiTfvHsHnHaf62Z+iiKXoUk/eC
HMcmRtNeQBGLkIHKEJcpgjSLIAn9ZiOe8ArkD72xUMkUFwWRmExz5ubUfjdkUnDTrY7TE48rI6EM
6HXOILTPcBVkjNuJHAl5dQCcjzuGoM9lyX1bSYUaKWDWkS2SD3LE6lcdxjpzuwGNVJoUr2iMRh5v
zt7IE+iLOUwRrMOjSRPrTuqyQt2jKMiBvkj53lOrG+oDIPPrKWTZ1zNGV/4gU3OdgCxlNOYZxk15
9jTS7VF48j6Jtz+C7NNJnxUex29itE9qpOAhGaYRuEyQxAOdOMfmLZdjfS9fjp8jPZX8BJtXUSzW
8gqWbgfnC5Dc5m2wlftP4z3d7qleUvmhBgxxPnPMFbrY6XSKggFfHzxHxyhBqzaGXVDV1VFPK3sO
xpoIQvS24AswNCpd/GRifF8taBrZ3fck3ExuwxWu2NhpzdP531MQsbJnlyc9nT3vzKY0d4vhusKr
DDsY0L84lAu5R+5W+DJ6FEJPUIJs+Cnqzbo/TChvcnDOk2Y9yMj9FXSyj63+mu/I6+/OYXB2mdxN
PGlN788604j5nzyZ9nXfCfbuKlMfNXI0gHzUoxe/j1BqaP2TWHH5r4H3EtMBzxp5NSs35NfYJ2sQ
vejuOG4a7Re/VvV+gmF5l9J25aetqHUPsseHCh2WzNOJ/DiD7gxFLQB6uxC3SwjJsCEGyTGdt2GP
L3hFaapZs2ONuqo5ZmeD6Axa50J4dmXYYfaFgVfkYnI9kdF4zinonGX6rzCazoqUC6lN48/e/RmE
ExqMmSqtKQgG+riDpQzFodioML2qgGHNMcdJ3Edxhbqcp/sG5LZcH9ZQdKYItd0uPhi1AcJr72Z5
5cjjnB6/t8iVCLgUqpzH/3NJ7QaA63fnPlUTYZ2169Jht8keq/DatdWnLaY+pLcPVacfffRyY7tX
3t9MMNUOfDzhHVyj1x6bZCrf1MExzGl1SvTF5eI/aJKDCYATCu1Rt4KyI4zWLcjzwdBFZ1xOPM0u
aRUH/JXI7VznEIYqzJ+yJpBgrYSGVHqeT4pUDnxa0WEe3ODP4M/t0mxZS0x6sT59z5V1tXGAs4Kc
9pGcC8Hy7DcTI+EMkPaVEmudpwRLCVUTI1eLC0QPlEbJfJx+SnBHoeoeI5eZDeP+hDhDtKY7KVrC
KdzkRJQkqDj+gjzeG+tmjCaXvx/3B0bmk5zcB7BNzQEZnde/iq5d+JYaFWEtdfo2OyNf4jl4KoqW
+p4WaqI3XjURI983EBQD8rcQXJDz9hZ43UeQjkZc1g4C6qMfTmeQjSJzJJTJflurmD4z0k5+NMHg
Tl5xNSqujCaC6cg/mdo3n9DiBEzhDBT8yhEt/RTHM9ia4FG0Jjs2GKkE0YAOVDAn3baTl66H3LD+
zzZlzjhAuSwmM31JRSauEmLplxeWqJv6Vy/c0ArZeoSppeMLUeSOndKtPT4ye+jee4cg7B2qK7Ua
B2FpQjqw03I8lhooEuRbX1I2qZcjAGKjatMynnyfi0DY4vf/dGazUXB0yywvRxIIN9qBsndVgQ43
8f/HNt8Mdmu/XGOdy2rsxpk0EJmFVYV+4UKUd3bPd9J/ot+ID45lrYhCyjX5+MrPzqMJAkUlnYhA
XBAPSOaMHAaeg9w1NNrHyJShbvFPAkLMNro6K8vq+EzrmxMqdtNWn110D3nxNLQl1gJnJ5o+jxyP
WzotZo6tzKasjPGba2Hro4AhB+Mmskipkn5q6xJ7BrrpjdAZQRqQEeyR/HISUNZ5Zz3OghSz7HJW
4rKk3DiTfEkdutHtgKeSaT/xCtEf316W+t6N04HAleVdt2qKPNiDxOCjw2LEJx40hM72yDIcZ8kp
qcwVlqCy8K9Jpyh8ibhA+0OP5vEgk4s6CFDe4FS1QAypQk8//5KQcIzHUGcLY/rJFwmRbF7UH0DA
i6MjbFirMXbYd8P94Mn94beGhlJraA/55qOQ8jzuQG5cq5Ptcy6SVb0XPrtTh4SLDuUkuTidmuAg
FpMibqyJF6czOC0wokjevfpOGAbHuPrWKnSdvzINuW0VISj7B9gKCr3UCjmt9yBXHF+np+k8QeDv
qr2QsLd9etlh0vxYm6tL1upjaoyFq8vQRIj7qjdj84puPAm6g3Nyz/1S9LL7pgHV1KGqp5WEIQQA
pKhPRe0ZLBAjkqa5ovJUMNoNfJHsdyr3md/N1RYXAfJ5nLmf9k4IYEUEIKZ1MvQFeAnZZF3/wnnj
kw5S8L13jmOLxlV8JR/0+PSWHd5+DFbuq4zBPx3lpY7+DPT4Hyw3+5vOuczsLrji5gpv7cG+Yi6U
TkSLEgsn/6nuuFkzt1RXRyhDrRyt4M+h6mVnM9Y8t76zQ3IXBswOLhGO/4xqy+v0wkudOR6nRyvE
RZfEhfDtvMXZYm1f/MvSgMC8c8PHLAl0+JJPZkQ9HMePrNEUJ5YNA2iN+uoxAvL3pKkMZe0B9ErD
Rezqz98D2oJzP0xtjaErNslBEBCeIABQP4VJ3M8waWubqGf+gkX+MHxH8cyjokjidKyvyetYZd4h
QTUr0LxNC4hxMeBlthCQRRcmRGxwWU0Yr8zIR+X+nFiAXMna+0JLOwIPQcHEiPpXcPyvaZRCtxf7
XjMbVYz27e94Tq/QGmjL9KuD5dZJdkBS7rowEKNgK2Ptk8zLq55HpdMdLNRXQuqj3dLaR7InsGbq
ajVPbaLcoyVNoLz7hXFlTuFXGz9BEVtLeLKnkf021Py6XLY1ZU/3rFzJlDdEiwYXJKzWzcxgvvef
RWxp1hsYIqbTAcnxPeUhFsCxEmgnY5Ljrmb5RLaWI0Icv+RwvAhChbyfYbj7men5G7GmksJsiU2c
jWZMLSIirBgdIjAEeKfNozIxdISf6sDdM4DPeW83y1OpmhqXUGJ75KExR94wkBby0ReI91roYXiS
yJYzSD5blvGiSWpg3iQYIVkJtbc9vFSUcm2c8PJho+1QT/gq3FQfFi1YFwsKkYPmgxSAiRvnmvNx
cYduzZJFsEAveiwg3p57rZRDl110mYUeUUjrbZ68Vv+ZJH3OO8XdlK3c0U61GC5OwkJOl8iwruoW
UZ4bB9bFssGPZLQWNVAtSGw/CWLdV1FlbxGU9TECdtjsD5iMI0VQDR/0Athr3PDYqeWWjONgngiq
MkmmbonHQxaUs3ssUlXqeuwS8XwsH+bSwaIYBNU9KHtQjum93gBOEkC65pUl8AZDJmWUfPHn8l2I
kBz8T5CVFudhDUPqCDJoxFy6Z41LvSzNrNM4GpPlgJwVL8+K/suwSWh4afOivABL/wbo2iH7Tg1P
nvIpAiuqDQy8OWtqrF+P+xNThhI/usSlK8WRmkW+cXJztAaM7Jx+5kHYqkTQYf10Z+SOMjrPHhd0
trCZHUuN3p6GZh7DtpPXgjBmyFk1XiyO5e+WDx+Yo4Ao5UnAnkcseXk7jxb7gJABmL/FFAmrsSHD
DUIyr1QF8lOV/Q8pVOgoyuUlu7khSfn+kkzwzCMBnrtmOPnwYoTEKbvW2g7ildcwCGROaFybHx9q
8XJ0ULqlTF31niNi7LdzSOQXxGDlc/U74bl4ZzcBZyaRUjaVhHkgaT4vtFRQyEX2Jrfynqm5skVF
IUIV9yvY8SqVL7BngckiIsw091a7nF3t6Wcd3YRr0U7Wcv4ZquA1eSqAeq25SF/iK9AuLQ+okBbe
pOU5XKrbOjY4Qm82CkBZ1wL2rh/dvMmS7EBCf/vbsiFnt6tY23rQkk4uyu6zRhPaplgdZW43/6kt
Ar6lhBZeM8SMnOvEaFT+HSj9Ah6q7g9TLOlNhkg43xkHH4TsT/YMcPivNMNEdh+tmOAtFR7oWfvS
JYhaF9Z8q9s5xddSTAGuZavi6/rSJb7Q7NwYOcDx3Yblkp2jOZXnxKFPRMB41Oanlznep358piIq
48C+84/XI/MluLfERDs/k3xihmk2lz3AUi+IlNxfaXMzDU+Sz1pIO4OuTe8MgXjI3zAuKcRGyQj4
j585KyNM4kN9GZ0I8uNIRZT2gGZumRqXFnNX9YD3MUOF21HsiYS460W9cOpznnd8n3ilXN9QpuW8
j97QD1XBFgjUpyZnbW1AmKqnGOLoSYkmr96Rdk6ZKKeW1K6GRDCWnW3+QfmFeqYz6LPC6wbb4VwB
fj00vNTsrPIWwR4aFLZ9gqK6mX7KQi3MIkY961ti6w1GMNhlLV6NBSncUS6pMZgkDKq86XsVM12C
31xfBab3ItXPHJ2s3/f9NslNxTzQUDbf8GjkYGmMHxBaLhZQS5PN31L0ORkbDAfqJkNfSvQqFLXx
fAks80CZVExjYcEQbZ4umzUIe1IBt54dFY45rA/P0Pi6LfwV6f4ETSFyET+TF/lexz4AJaE48zwj
dsbhJ4I6Er+HPGqEwALDKDxPxD1XRACT9fKXLb8vJeYj275DiYHeJuPtDQC4O0CQGNWrUUTJ/tYQ
oBfvI8XGhlEr4deE95x3IbZrCjBCZscLgzNevYU+m1926WsadypvtYvhFJ6xofhWBv5EZu8Kgopq
9KqPZ62+3TCaoLJR3f/yR+Zdy43/shccOx4NQzN0BNevnmJ9N7grrQ+QxrOLryYMi6JCunor+R8W
F0FW+vLrDrnGwkK3tPV33gwzAtggFl1dwdE9sP3tmFnfuYnEcEps6abzwpXUP87bdmmV8CdaobqK
4p3rWMLawJhoC0oz6rR+Cob81J9aEa1njEYISPdrz3y87gEdXLPnkZqfidwSqXDGcYDFHMCXmbne
vOetxWJjtedOnqFnswbxFRWpwNSV7l7vHSpu3o7dWtbB2SPvW/NfZXdtJvq67P2Uc9gnS3tkP0nh
CmH7NONHuTsKPqczbBgI2YfvAJO7rOZlf84n8RTTfr1UaYajWLfUqntn2dgO2WkuQduhsLOmZJeZ
mtnPuUiJbHCznDSa4lenhavVBcGXIWJlugqERlkNXkoqdf/24iWrQkR4Gsoq5KW7jM+I9tLVv6Bl
EeRYKG75MdUXXAz3KQsw/3D44kGgBvGOrndBH7ve+iGGvT7Tq93s2iDdd6ImiTh+YCgWEfIXAL3G
WIPxn6tyeev39ld1P1WwuoDJhsF4Fn5cGB5r7tFNvXkW/XlksKjoaq13xpeaaqO5bYT9js6EMTz+
ChyzfZ0JZ5e0xKpC2XnHcO2plVw42oU1CcDPUvm9WZkd2K688q3sWpFq5BEcrg9WyTUp8+lD6hns
e7ElCrohLHMA40j4eUZ7ZSx4T4K7mgk83O4ugnzpBK9B4H0KvgD/6lD5DBwVPko8VplstdxONErs
CyywkqmIuQTQkxXUvVvy2qRozAh9VhBTV58f7JCcb3BTrdpkcGj2d3zMxMHnZ9VKm5Oe7Elby/Ya
l+xdNfai/+4MAznUbFTvwND4J5xnRaiTMo4XS/jcrhkvCGLGcwo69pGBUt7QedttgMoAWVzOdUnh
SuEG2BjnYiR2+IMnAgoVwifybuGQSkVx520nECb1FvAfd0DvkEJmtSila1PnkHnbdXtMFPBh8DVr
UJh56h2ar05jmCYczIodBbrCQsflYtoCS/8V3yKagPn5zuxhDnn4mUcrGozVDp3hAqhcKq3cjXCi
I9Fa6qm1xwPk40FPpbI+goZipbEciXwJWPMS+Vm33KclErA/28I0beKrsaB2Qm+swHuFeJHcLwRF
833kHQnh1XIXCjL/+GXO228b6yM8H7HRkhSmG1k8ctLhZjfoDaU/0rIOG3QtBN6VxlX6zUynmIWW
t5LLSz14PzLzx45KWLrjg4K4NiS45Og6O/jE8nCb5PUZZhbXBISWIVDqqo1oq0mAfBj3mgFQaTMb
a4wKhYb4b63SeyfVKLa4IhhqVfghQBK9DVjb9ld6GHnCXMoLYvvwJ69CmKJV1/gVdBJJSdJE1F5z
/5/adgqnjEoCnX1KM+P5no+3wlK+PcKpCWahp6vc26dBTT+66XcZLXTcZCsYSQ92Zb2u7PW/5z4U
PpZzDNc0naYdwuz1hPYY+YN7I/PMGjqq1Lxltek0bPAW96a2mZeZiwRoqRsloPRGTM8Zmqrbvfc7
pdRTl6k70P7iZILMkM8wLuQUmjP7ASBFTtWheFKHGOgdH/4HgPcBKWu5rVKVmM5rDdNqoe4r4fap
NIJtaA4VWLZlWPyzcvLSCeDnSYmqYGV3QlCyJbgANUWDRVGg3riPAsP9KZ4KryEhlQJn0Bzkuk/C
E4y+cRDkocSpdoDvKl8tK+XJmW1lXE5K8LkDbFEqly0ES/IUNm6Tehd502tC1xtDPUGVFOCiU0qJ
heDM5+RLW2/fi8jwjKEzqTZ+h/EFmXVf82z8PxaY706g2hvBBYFVBMlZxUEGn3Lv/Yt4E7JIobhJ
G29V3b4KI9IugKrlYr5/xmGmDkTgCAcES6BqN2b6DEA8Wf7Rd0MyXZEQtWDxDCiRQNuaaegu9xtt
BmW2CFrcnBLyknwEw88Xe+YArb/XPt3JtPCmX+8L9x49UYex8M4GiETFs37hdc7nifATCypBv7+s
JVOxMAHP0n4Im7ioyule9mGEwwaxiG8tuT/z2+2qANKE/QH/HOjka0HGgWG0FE52qmKF4WeGs7gt
tj9oEsLTuKfK/9D+F5lVXlPBM0NcduyDpxBc+Vx6TFxNHLbaJt29xu2GKgb8o8u32KcwUEv+YxD1
1H9A+ZfSS5e9vWoCt4iIQxyq1U4BoFphT+/3g5f0lyBU+r4t4dzcwse3+2/5piUmXdOKoAaFx3Ni
nRpTqo2SR4A//qZKU4z4IAKhaCHtsgYdY5V6jOtUY2478VhVrlyWFixg1xHb0UTMkZZK2myud2Cu
9ZMLV9Ow0StV+dm4JuOqSjCFVcul/zcTtybBs3HAxAl36XM9PwBMZZvcCXE7FSyJObc7MDm6EoSm
+tU6HodP+mifBIxlADZ5HZA48DN+fSZ7HKhQOPvsZFnkjCrDNkIFWMtEodV/dDQCqwTZ3F9HYk+m
9n/8bLgsCG8JJ8zmCG6KjgcUUzO03NxGqz4Ai1o+8UTXrVGEy7cdiC5ug61UubZQUdd/H0BYJX4n
hagDIaxT1OjZ/Q1en0l9MaFg22HVPxJq4357CoRN+XfO4YXfIGMd/E9gDJnjX51/vdlCX93HKLSZ
bwlpoYtgJjJgZhhsgYn7haiACV0LN9/zBX65/dgIa/Htx4zk5u8sELq3XX0soiYIsO+iHmljT+VQ
ywVjq3v1KsTtE6mISpW+8FvDLzMzgX+MfMGXZ3Od+BkfGCT7CZSn+pn6FZjyffaA0FKwfPkbhTTK
6antTqTQLMDyDkTIBQVjKcEHqtlK50RgUSDKjzY+ZvoNw75mXB0qbUq51FRCt87RcEhBustghW+B
rDiSi90i8xDZav9p5uJW2GcJ+YHeDfWGIfL0BJcFV4mDwpEsN1E/GlCml8HdYhqNWXyNdZOZRzMG
2wk2VgICi4Feh40VeyfhCZKRWMABD+IEKoC58G9wT2af307HK6JCJKTL2GdKW5Avu03/BLkw3/oW
dA+dZpM18JLODv8esCuBmONHQtHU/tuBOExCCp7kGJxbOknjKbisl+uKl96Pzmmiyjpn2qmEBK1M
UJU4gc8+h/Hs3C4GjD8mlcUllcP3R0b3RbtHoDPDD4UT+ahH2ecSTEooQoch9/mRUTz33VKL4HnV
uLO49LGQDgpS+cveqizkuVQSrLl12H0E33UyJ/Q7PznNril3314xD6Hhl349V3Bt++lhZnazPQ5g
gcFn/SyurpZ/rr3VsL4k8dAOCQvb7FH5rRoFehKaK3sx8LCpaL9Ehxkr+864wEnCo9fY/QRwQOGT
jDhZ3fxjgI0Ivt4Hlc/rMCudpHJFCwlvqA6NPjbXg6IfsVtFJDGSaej7F/zk/KQjfgv6QstlU/OZ
lXp1FV5QAAFaSU8kUs4BTX2BZVTkNPNWu43cA2k4O78hn2bLzZ/NM+o++E8nbxu6xdFtjXpu8C1J
0VPXOSvE7pYV2PbamrcaXqpStl5ZmIl7kpV3C/lGAIjNB6EKS0JD31rZHZf1QRQSzxDw+FPHwfVY
qSzJd7lrkcWYS5nTktQhV2//4ihEwEEhX2Y80g01jH6FjXZWnKpIIHNfnmSwqmX4pWkO19n1n+9C
T3ws7JQYUIThEQ4IwH0PhaYJLeJqUQJe57yzh6j275Jdz7fRztfzvNJ9lk9tJHmSUzvXnarRY3wH
YE4YIViE+yVY/xMfb5j9GVuaGFNajVNno5S081GSrrRuyDcdQYAGjDsyOz3MWgdZRVCa7ByygfW7
ZbpRgvIQvnjUU8mZBnWmamUoVHd/BDwYTIbIJEZa2kDFmrxglCvsSMf7wfpRAMbkS89341c+SY8v
yo6R2aVqgPPhXuEZNEPuwWUQowswLJdyfbQhwb2R0h8mPLdNRjd4Oe1bZ7xhvloaKPahSsjg65FM
xCwtIT2hBuLtacIzsJQt5FYWtvQv+EwlXmHzaja/FcOgjg3b6ZpDhCNE1gyzuqjwxFC0Fz2VDoNs
0qmiGxgylu+olglRNqSBjBX+cbPHeq3YiW530cReY4hPdkqSRSyuQdZFbSoKyjS5Fyp8vSf4GYhs
3Da9JAF6UFR38R3XxI3L8r7yBeGlkxPdJk6J4hgQlRMzkgJLDfPiYUrzuz5Zd4w5hFOUOECGV0Q8
J4i8vprfDED+xOEQgi4X330Rf+CqmdtbeNyekhKqqpL8JBd8NxVTxhev0M26HuSBFr56Cr16alTV
b4OaufK2r9CZRJZiNTN/+9Dw2uMQO5HP2nvMBFm25favzDXTpX0kynqZgSEhfk1nYMjO3O3f77l7
aSJO55gzCmvRm+mMcpROdNQUqttP+eUtHEJAyFM1oEzmo0+IKICSP5VXcZaEtWZWz+3HA/Hxgry1
O+btaqvcKhpqfGbqDAaeB+OALYxkxXlPJdtGvFTnp3iaiZEpxZ9IJGVzHiBWjmku0bFph0vyjJ6v
+N41Ga2LEiyMMkgeaFXK1+NwXhbsT6RAftAMU1D4h7UfY4b4/8gsQumyngaOXC7xzGnHeMxo3fGb
1MS8FK6hCBV4V6yg/VbJX5DTB2hmzRNlomwcvTJN1iIiUV6xLHISzdpizUZNKEe4MVXj63fRWwJ3
MqD0Yb3ayYnZ5tUQwPNgDHVGamR9hPfuOSNybtrb8UlRDfdVIzUlJBpfGnYCYd3hjCoBHhn9UGoP
0Wwr7hiZjWTnAOARWlPrChZQjT3oyGRgICDrvzk+j2oXcLSYyILJLeTaP+sqmktKvxkH246SW/50
G/UDRvpojclrnq70sbAMZr4Ktrg4JMTjKJY5lDQCs7d5MmgYXH89lKsZq4236OB85o3drNdPSClQ
5F2BvQ3wC/kKZA8OI6QcpzGF1TUlH8Y5TajR7MioUyURs+mC7UVVVeiz7KYXMc+WTrn6H0ekyaOp
WSsdvh3qOxmCAjsCcf4HMKPHqKHMwI+YuuQ7mV19zhZy/2dtuDqJFZ63LIct5K4bn0/V8lvQ/YPH
3x3vNoh6rrcmsUuIchas+dZxfoZx96AMHikWhvtvqs5vOu6XF+AEhBf3zTIQUcfTxDnLspVyHDaz
lpM5cSQNiO8vrNaWPdYABusmzWZjU4Z1uue3KbgLhewBoCF0BWAk0f4LAyw1o9bMHUCT75CFweRQ
LsyEb2WS7Q0lR7moEnIhyJyrmM0G7XO7o75UEqPnk2G7tjRAAX3w9sgTQfGUYsLG/1E1JV/56dsp
12Gtcl2FgJjifpDh5+N7a7dPnZ60HMvV356slyhQppteiFGBr80SN/UzgDLWAE7H1NJ9GZY2YwMc
QvsxaK7+L9ydUGQR2lvJKLOOCaAcCVA9RdRmHLG6AB7Wngi6OJJ2jZv9o3/svdqZ6I9cQSrnPpMg
3+lnOgKa6OcgrxklA9sjM0Fr4caNe4yukZ+Qi4o2W6gy7tD+Zfab1JuYKYckjeSBEIOKIyR/qSvM
8xE+LduZhUS42x+MkAlmzjoBCpbaHGW5O+RnJvhb0lhwaO/DPfvRDdeYA3tIw5hosGLXpvExzdNU
BlQkIflgjW5SWwLG7+kIFLQKrKWkCskp1FrvPzHdkYEYzuo2swcVoON2+ZedkwdI8spdBxOzBoNe
E8bbKW3h1BP/U3B4M1mKaJYh/LqiptpOcMlueC0rDlMrjoa/g6NrapfRgXbpWnH8v3Y8K9wSCMcB
TqVU7Jo4vo4ZGkphxZqqSpFPC0B0+5T7CrbF2A18b14ONwWFCdnFe2zjYnHviIjvdQLryY3cSdHu
0VNaEQQYMsD+dmLwu6xANfDtNXyqTqyAm+laNmbXgRBHwHH06aNYCp7ea2ONkncVEbCJqkJgKcMY
/+Cf5QsBzk0qWuOSLudSetegZtfI12LUpk2WnlETUlAIRAeiV6RCgBrpre0L4loZ+iGDRsqOCDM3
ak2gL+7PvyJxReQr9gYR+C6xnV6ng+xQQJ+Qq56tpnG3Xq4NJPh3mJmp67MHsQ4V0tnKT6fxW6jQ
K89PmLrriWave9m/JAc+4A343PrNh59OFPaFtgUk+tguY8MluN1Zf1nURTSghk4nbNrmKq3fr357
Va3EqDKH2I6sRPbiwaa70dnMiAI1xmIl0fuKbONm9dJiZ7QJ8j7a3BG33g1qO9z+wRXFW0DnLTP+
ZaK/I4z7Ww4xFMHQl2ajonNhcVxGCmekYJMlldQ2gG9qTDO0rtmRKWDH9QCbRanUDLpVBwnrObp8
iJc0xiD17sQDUxnpmd+OVm1dwqYSXEq+ARMlnbDnoHfBPj/jBbeGXZ2k4MzwdgoyFUIZ+QujDF/A
8/5Xt1gcPCHKxMgWGgj7crcBoPu3944VqYez4xaF1WpCUXCovhGGCo5vLntrmiypCzAoKTBPOGtN
PEqSZ+mFayU/Pl0XO9hKmXLKGSZdAB6n2q7dhD9UtoeX7KLiROiSb3Jz/sFq72X3+5Q9rqYhsX9K
M1hvA+IBlxPgstECWFbZxKQlVF9JKNOYOD8cEYpCNEmzw9OujZzs6AT+/+XHWuRw1TE72VG4K7hs
9jlciOVp3/8viHPl/5j9LH2VGc2eYO0Ua7zg/s7GkCxVQ+Sn31tPMRS5oIsCFjS4mS8q4qmXW1PV
/ecrO8LXzAGY4yVaqOUWKNpTBL/XegXC3KjK4lOYVw/Pt5NHxLNsSSgLR2bEsV0jPXsUUlYSDzij
d/wguyqScBdxAE3xclAiDPyWRScFJ4lHYdR/zJcTfjTvZzXV9GxLYEYjPVmZxCBxH/zgInQTsV6y
+jA1VuEQb522NtNS2MLf5WjXgkqMYFhalX25NL1y5HWpi3RnjVUtzMA4Fms/gwqUSSA/BAPtQXfE
5/aSWykLmhvCJMUbxDKDkBD2D/+/ms+wD4EvpOKL47Gh4GAI22nbHUIh/D8WYH3nj8yJg0AV+yjE
9kDMBYMmCisZ57KKzNV8l9yTGvDhYkCup6hle+IZAoulgIkeIej5TQc70W1bPS4z/dIxlck6EJMf
+T4+izN2hua8lmDj+yzkP3XP3Su4t/Gf35C6GXFi2wK7Zk6jdTNPN3qRRTuWYbITytj48Hu2Z9/Q
2O+Q/QZftwCoyS5qT2h4gYICgsU73JdM1G8ykNtzy+fCdce9rXCOcYTJe5Ef/cKmB3+oMT+BBGkQ
HNWACSnzfFcP0tWKKrUPh+5RWL1fPzlD3JKOMxZCL1wThbwL2PGBBuOnCclFvBcfx9GOg5O5Zoyd
A7vW4Jn4Si3zzKK83zKqYLAY2RH9601dUfMKfYO2g31EoqIxsmA9Hv8xkcH0Gd1LPcbLRisHg4Jf
NAV0iXiFaBMG6yLKdFwLRlbULiKWoqkG3IUNjsmLSaopHUioCB58h9XVe6oh+UUYtI9y1oDf2qxk
D5GOgB177W6G9SSCSsdioNq+Y7hD2gn5eOIH4Gd53DRgqDZUkY8tq3TkFZYyBYB9GbsoUxhg+Foi
DO0uawatMCemaV6i30YwMWNOLPw1Nv9vQXheWFGlN16ecsPczR75RS82Ax4yDqkfjOA9Gm7yrqmx
4AoUR9sOWNWBjVpaJDnSzeoEL0oQXmvC+pBSEjM8jM7Xd4L+tmFDasH1IjbVitqRJk4xpcJtBCJQ
bFybL8WhG/RA/I+CqSwAKWyRcSKZ7gCdgJgqLZQcDk9fwz2cIAfQumuWf1I00Lv7tzFRmVEcYvgo
qD9mf65M2aeYhh5R3eozd43o+8mxeHwdjXVsMwEzVzDSwC0ppbgfHZkiuxKqsqlzrPIS+IH1qs86
Xj4Acay/+RKT4bm/2R1F+v9RGpc0af+WZVbXbgafZvfN1/13IPqwxaTzLPFsBf2F+/oP/pnr3NRO
Pwy49OJ/2m5HHXvroLbYWbVDFi7qPfg4hEsGNJ1ojSK7Wi3fW3WDggxp9SkikPt/jeyVrLF9IPGu
4kGaNjBlJHgOVSXwyscYRYxTmEc0BIgWcFx667/Im8PtOwXjjzaFaXJnUCQXdb6Zr0ZV/+n4xp4n
xG7WmR5yJfINGhRaLucLHCB/0k5weCNG+4OdcwyxDoVEvNTeF1XlGYuiovcvNQfcc2t3hfYiXOsy
FTdlncVNTlJKhMPv6Fdg2+RWGWUEHrkcNOSdVnmnARzu61eNJw5blpSrePo73KcC3EYObfSNK9xW
s85iOeazH30ePkAxDPnbcJ1IBk+QVSwnXO94ZL5AztCpFpqNpVZkvPEu1gDJ35cADhBiGusqe0Bt
Sq84Zeav4jAE24pSPljxnejp2E7KIEkBxQJOWhOdPAD/iq0tDiJTnClxJGCzpZAtsskSLidTSBdi
ZCiN7IrYxcm3liQdUd5gpIG32HFCxaJ6T5XULQR0VtWwaC017j098E9ionqtQDCJRZHclqaECb9E
X+cQbeHnlb3ykpDEn8Zq+DekeRAlMJ06hsnufWdU8SxXqY23MFPieML61sC8NwHulin0OYknc1AN
Y8ip5v8Umb4+la+TxvZu0Qdi4wu5osjMvavvAaTw+mA2NVt1yf7pcpm7EosHqxW8B/kQNQsGkUiA
ckgb9D7L9uC8PbHC3jVbGXosBqly5i1ND1Ztu4nmWOyUDpOG/PvBsd0Ieuj7uCuc8JHSFJiRQdgU
e7nOfc9VNSWv60Buwv0VrHHS1m+N/k5mqgPtEmJVF3oERgxxmR0P9yBvKMymOJe1f2PTBqf9Qp0h
BOE4+kmBCMdGQ96tX8yME9AIfZj5wpqHiMPVz9k53PGlHGKQQcYuFqyeBGnZoKKWi0RHXDK8UIeQ
hDVBNaJRop/h+V3r0WPXoUmi1c+3zmu3rC0yW0CDKhGShsaob1Jdq31ZJwwj3u94zbRCT3BavyvH
pANlbLjCwf1nrv033Df4W5Emy+lwy8lzmUbJccxj0pgrOqjRsqSc0ijmP2/+ocyXFXSQF8lRCFQo
lTQNO+UgogBlrg5NqoiJmNH3bO+6ypWh5Afr3yS2cChBj/xQ4O2HtQsHjJQlPfc/pYf+/g5nkPNj
V4qVzW3tJ/fre8dH2+yohQOkvR5s1yCjfgLIfc8I++TKLfN/yMt7P3qqZAbsKSpPd0LVo+2sL5z6
DJpqwjWnz8hc8pw7kJZCS8sArnvBxVn64oJyp4KZv3WrrlK8fkuEP0sEEp4kUlpKQHT6ivN3KAhV
cwAWF2+qyYBjmg8QERjc21PrR5oYxq6owDm6onxGvlJD824rd2HJ3bcqTx7XF68Uc0Xw+AemUEKX
ewomuS2x4mSrIkbwdbPiYSAqLal/iKCLn/tmnl4IgDbX1b/z8/ovdnBf5MUXdYZGMyGep05Jqxsb
dgngAF7eo1GFCzzDLsHIBiGuMfCusvOIFBKKgIJgUdSbWD63tHRPylews2aHrShK9FKLBsEgwujU
reW1ayiQJ4z1pwZ+gtPMQWP20yu3LdSwwhrx+bD6rGlBWG1ejFD2S3l/1rkuRC+63QYJ3cV0r3gg
OZIfxL87PuYQ1+qDYaYFy08mASb70Sl5jFGkmx8OJe6NfXGTC0d3rzHKk6eK93PVGK0yMT7VMUN0
XPNm6li7rgoGAOXHO1xvhgYWF0GPsBlmloHQXoyui8Wpsn8e5h7/sqMhbrRcnXUQdyfiGyoZfbPu
/QHbl7D/KB4wxayTNVpuCaq/oLAj/hZZAUXZfXMgz5VyQimfouqLdvFj+/teVyuT5znJhT4wePWV
5SXcK1hOPnlVq5zAwwQ0x8+Qq3bNLY6GHNIXZy9QrwSl4+CXrDu01xJz1L4nIx8mUa5xvxHwS6g/
QC8ZIr8T5yDMEZqToR/BesjPBMUo50ZgIxesbzB5UbSdN0Sc36Q5IJwkVOORmf/5YXktpwNz825i
WVUH487wRR+++IX5KM+OTnH2E5+y9PbxHiLTjCa2iOxdFlIlgkyTryZ6/0zaV0Zi3IpFk1H2XBlt
aUBCBXVLhf3zUDoApzuAZtPgdobCrdHnTrcfKtelB/szeTfjkmyCCcOq+3HaVGsr3imPt7qUrPn4
ee6nTBDy5zhbE3VmDXNhySHhYnWKgzig5Xsgy+QyLMJtnI1WXo2PVtDOApHEfCYmld0vKVxB/Jlm
W40Y1q1H//hAvM8FpvvV/qqxnc4jWlqkc4U/qqpkh/L4ByLaAEuGI6beP7mL0mALHMMKDrwIGywc
tYA/cs2AdAjBiPCxfbCvDUyiocmEgPDn7/nTbZzu89uRaJO6BRgYmJffLMj1jqAGJzurcaa8Z1Og
x+L/gGYTIbK6roxBroqvhbD4Oa+8b15B0TrjUj3XVRuLCwDvGS+R6XuHDVi8qIZ3NjvBMBchPo3F
E2SPqEcTMVur1kVKA6u/4ML7Q9R5jDpNh7yBS1j/AloGWRBG3tvUytkIFXlyj2xsRF1qSMOmM/uT
sVjpYd75aMMDMAXBWFcAA02vSq6pKvhg0pFC3Lzh+jlyUk+6aZTGHQtlB+yOZVkTMUlCfkkYFku/
Ae1VRC3QXfJJR8aJuCmeF6FhdzKR9o/n9jgV0QqP2U4PLHQcE3arAKubFIP85ArHNfmAlfRMM68c
8qR5dbM+wyzo0ZPFCid4pVLwzrWJJPu3wnfJrmzBaeY2or7RML0z9uMkU5kHBmZA537ekg/CyjnT
w/un0Bo2GLcHNS4OP3lPjERPY4y9UQxG+5q84J5kwqh+LuNkLhF18HjJ9tnQTAS7TJanoEwIqqnI
peOUHrLpnIOTrDRKs/Vertbm3DjmBQczUzfiYOlo7MsEhlJb5xOLg45Bpubn+xFU7+WRnNsVPtyH
AvKqGRaWlU9hFlxEZ/aMear6r0sXRiIXV44dXdv+IbcHp0SvnL+BfVNsP3iiVtzDRUIoKertLlI6
uf44Ss8tJJcdY4SkIj0odZdZAvMk/odVHOtXzMgEAkEDtGI8zXV8EHEeT2/qpeJbBz4//kvN9VYF
+7TD6vgtD/+AuQrAAX/WrShx2BPeXxicOOAeH9LKu0PRFn4VoTpXIyqpDBCuj9zawjuAJgk1FOfo
fK+lvJ+71VvIz+AMOPg1k8Y2+RIDkB4IuZBfB0PP0SzWEQNNxdYGRUeJJYVwwUGctKNWmsbqgK57
CTicvpI3mG3B2lbl+eHt0YfqzvD4zV9d+l6dY0g8qnraR/JTbzuUP4cGWFptlxFhNnN2WdtL5eUI
Ep3lDbfwF663KcW3nmPkf+ki8elTvZ+Sgk37escCTWpbB9vX9BWvGa64L9UM866+opQSmdz31h/+
90W499Uvm3f/2BjJFOMy1Xs7Ox1lFZEWoGVQ0ypVOakIg5CJbuIlhSfxDxoUHmCNt7KVniNgjsOf
04ABe6rqUseWc95poYmIbA+XgNEHurUE6i+OLGlAP9z0kOf4VhLB2FeBN/PGkjNLbDtxMACv7XXW
HSi5VGS1uNZwgNHzhYFPcJHnlTUc0IWPtiPA0y60HiBb4Xl2DqEKI6d9vssZTRBtJs+Zf9Fq348D
ZkZkwWfMVzLXDDLLF1lgRVrvZnfEoz+hAAmFpiMkJbV3gwXlxlcvZU6qiCB5dnVTHctxS2FnZKlJ
BO66VWqzBPAO4ln8f3gLaL3yeWaIe+m2J6tzthle3mgCRhff76Bd/nTtcCwqN4wY1lpK5+EqD6V3
LmEtZDut3PLsEa2nzJI07W0tNX/Xn5s3NOIz3HkqPdRbb34dQOxQ9EcZXUj8HIXt/FD/l/5vzX5S
DoB0G0yQXmnqN06Y+D/ryRM/4J1V9kMggdmMgUEwAw7g1eFXutglJVjueRjbZHR4qIHPdtBhSSan
Fz+Ckvc1l5dgCpT5FXXT40dxKQKRuT/wEzWTxVLkHeVCrLw6DQ+sJL+1y3zBac9WUhG78WWmrsTI
+Wm8fR8bjLder4M+8HkGYxR1A26tG9Lmv3ZfJdhN8uGIgFul3hVqh7USOibjmoLXYenvQuwjwbwA
RfW8iyohpqg+/dubeqq2738V9rT9yXsHBSiEKETKgCDx++UdjTukSc1Ili8Qwjs4KC/1TDILUORU
Egqp0pDByxjeNLgR4QJyqD3tNlDYwz3irQiCeSeRXNa3/P8tqeSF5kC7CjHvCR2IkAq/+RbumOey
S4pFaGzb+jy3DXz7ikdaUkJ3ljX9l34hFoECuhIEIDmxSMcrWK2+/IxfSi9t1+Id+jBzCCp9pUWR
uySRmrnYd0c9FJaU7EUb4Wvs4gdToful7seOF/c+9pL4MTURzIB4Rpongi3lxm0CeXk84pTRN7iV
+BUwQL2O68nkFt0N6MoEoaD4JfcINC9kcg3xEWqx+hps0OanXqHBtVHLQRraIP2AA+1ZH19Rdy27
heOmzBhvh0RRQKGdsE+PdOUtt1YgntoooagvE1o3tQtdwPKe4gBeFv7uAwD4vQUdezVQhfBwU5aG
K+8vJk3iYxACMdPlDXkPUaY7qnJ9eZ8+hG915AZtbaDHC8RM2CDxOEcB8qNNjgMwLyh/US/qtJ5B
K22OKWXX1uYC1vWH6wEMTZQjWrH7VzKYkCOYdn6+fzept5sONre8zAiG2qVi/BY2CIaWmOosrv7A
0c8C1nJOxBZgBFEgvxbpiHKyFahnM3bErW38xxaAcOv8EuHf6dSV0IDmOpmSSthKJrP88ZpgnO0+
WQDL76fSwmCH0h+RCkL2n8jSC9SjOGCTDGnfXPcd+9AyQQuIBNuVXg4KGahIGSAtfIDYoGq34K6t
hBrPk5BjFjayQmIifPxlDswlyke47FMX4uRbii8+dUIQXEaT2FIihMAMdbGkQwMMhyVJ8zy4AxbZ
9mgM7AZ2ftt2vYUG9ZB7dH8gZC6J+zUnIZtgz9Dj4uJpEs0AyFIeU9aacZ4LjYjHckQLd9QuXTVz
sKwLB3l57mx3TOuTBA+06IcEPAOT4FP+79HindrYygfGzLJhblI9rwTQNKcIiUA3/QFYem/1ZX7a
DZXAm+LGMzQ5GNpvz4dR95TxGU9DInBq4dqhWuZewKy1Fghaiwf4HTmINKS5EALpU/lsxs9DRa6I
wNOhQSCU1PhK1hhl0pshYAICPUff7AI7618JT1eNRCEbAa1MEtpwmGKie73K1XK7ADRbjUdU3MlB
Asyy4QXHofc/N868Y+eDgtHRn3lqbhoe6D2ectj7W6SCkc2FnHh5hQL1P5fo2a3BxgGPbVtdAd/Q
fhOvOP5KyUs5VaDTk4HJDtrZHtfpQQHWTgjOxbhj9r0rUDpXTh0Ta0hBnG6sS/9S88yfFyIJvDkQ
bNUv4cqGCYdqga9lBr7xYTStyy/ncxB5mrfVYoLekZ18w+s0lqr00jk/JixJgeG+8pSZTT+c/qIf
m0EfkhWtOk46y80SJquLOOzXOVE+xuRvMio61CFnC0E/nN0r+og3oDi3OpFOJDIaPsRPk+fRuNpg
DBl+1i9AGe4nZ7pA9iawfJ5vHbSogmAEiQhQ74s3HhkIxaSY+91I/UlEgcYo8MW0ns51V1R00w8C
J6Srz+rfSVnSC6u8CgedtY4NMoHP2Hkb74JZVSdA6mZ+FMeRdJMDYFj9avcyxMeq9LKj5woWP6Ys
TgdAKOPBsCB9KJ6Oy+GiA0/VpH53v+MrCsPOb9ccJXtJncSuAe5bi/nf8cW5kq5c7gNaUsAGE1SG
jg2a1YT4hdwaZEVGCEuN4/jE7SB4ZkxsJLwzr62XWcSWvNod6JJc2Imz9UOmfQwuMyZ87f97JvIB
/tYiiVNBKE8s53CTNr4ocbvybqeRSA8KIYTAnRZ1xKfhQlfuAq5fMj0RByrsbT8lIkx1/SIvmAKH
QGlx+q0pr33wK7AW+QWDwpVg3UQgraWBmLOFosKogw+iakBuNFNlEO6F2qVdHcbEkVLHNzbdu1If
PUK9k+lO1Up+X6v038nLGUMpOBELA3rByHV2tCS7DdfL3OiD69ydO91nkucnI7cyum4haqKiexH5
7wJZ+XqYny+6OGJQ0Hs+R5e2Q7yYCDDJxnVG01bU983gaYQxg+Tdu4v91GBoplPlTNwvrOhj6t9Y
wKDvovG3z2qvd0EQTN6rzQm1TIJKAI7IEJsm3beA7KvNHUXCnHTcel8sUBNQy76wuSloeL5IDgdE
dEHS987txl5OcDKMJ3EoB3Qy3sbfAZy5PLdmd1CYaV/bK9hfLsE+/wJTsfx0DJqOocwa2ERA1L+L
4unFyZNGXtOUdQZOXp1SWMaWifr6Be9xS2HPO5COqAF8uhwlvXKMqCfV1TtOY3/jYxTfQoBoleAD
XAYMq8oUg2k8vDVDax8/TIopi9PkI7wlnFG5VVHpQFZwzSS2/SGrTEUXg/P5EV+BloUPyQZ2BMNk
ltx2qMF2HqYTYrggfNKCKC2gTUmzaMEFKiZIJdvyBUMiQixbNVQirmnIrEXe0HRxkCHtTkCfDIfU
vsTLaniyRnNSMN1XptSE9M8VWS2+XXx7yymwTJs+863bK8BOXm03D7U5ZScybLPebO7StauZPQv8
UMuS4fDTd7nDr4y12yf9/on4PR4/odzmFwFUe7jh3gNJF/4+4M7qjpBzCPq8N4O8rMWmKON/0bgP
npqHimbb5F8dAMUulayjkG+m1AcoZ8i+ZM42N+nC3XwzN2Dg3thqa4mzB5VZ1Ov7KSOsUS6JyzwH
6Zm+Kw/rdEkJweMN0Y+po7qBcz3sexQuiFMRoI5hPMaUd6ZqFpkLQrlJ2jPzovIAtK4YwHR/I1zZ
wWCBPUNsZ0dOYH8Ov6iKZrPJZ6bOwB1A6RG6ZeDpile+QD5j5XKsjravZSg2BQyrWcUICv7BybGB
jRUckIuUOqUHeQQBbUmW9iCQzUr+sRCVRSwVMr1hp9pMj5gdJ4Ipqa7ViAXRVRJXK53ddudrOEat
G5NnM65zLG9XvUtEmc3c6Pz67Pehi/aOxpMYH06x/obDwCm509YM/DpIjfefZuFojt2Kt83fgRtY
pGMiqw9sMoNhBqt+U8ajjr9+vniTfr9AGoVr1//QvLSsFlkQP+UgIm9TAf8eLNDVu+aqWRDtLNie
EPfgIf1wZfmHeFRDBy0i4uFjEq/sUZjwC6DZmNoUOlE2GuY6x951oZ2mVziUaZ7ZUj5VsRjJiwls
D+MqB48+qDW/4zDanmIKb/m07SM6Xb+EZELBwYIbH7An6pfD815CjueR//p26wivHCrbkpEbEykC
4T9UmCoktzx+FRThhqMu/KxLQe+wAm7AhElP/aaKw+C42fnLyh+eTbl5g7YYVDvw9Mf7MpzuMjI6
ZIuGuoG0/uSTIebLimH3YjnWJUvpmVhuEK28stlxGRCuc5bkdrT9zmbexqhFJsmN4hmdE9gCumlx
vQdrZhS1b+OGx01uisKAtBNZMjPtetB1XvYy8pY/Gkz6MP0Kj9RQKcSYhBN3zj/M/0oDwpq3BnZU
d/f37OeZlA+U1cmhX2JYzl0T8tXN9cfNHD+zYZGkxoOUp2qkR+OngpKzI7R9BSfKuVL15vluAtMt
JvHTaotdfTr1ypzb+49DWkpCqBgpEU9EuB/1J9HuYXxEHAlFu1CcII5s87h7TIlMc6b9O4vWgT2B
Bkcj8ifHNotjILushjuJdAFme7BMDVmkmuexc4XaCqPvu/ZmRtcsyFnAtT6I7okeMajuzaQ/nl8Z
i2sjqj8BU5l8yI+kyMFfPCcWsAfNeQyTVdQuwWVEzPLqdw8+BWPHS6LLLggY9oufqHvd1NdfP9wv
2mtXvK8R34+MGfo4GTMvMbFczcDaVXp4LhOOEw89Amu2u44+ABvcuQ/EIw/+i/dIINhgVnjDn1uc
ozUY8M9zbooNrVL0dsbZejIy0RdYv5RVH/SWsS4uQdiLc7Z8zLk3NtP3C8D2v4y3flWzyT8eumdV
S5qns4NP7t6KVG4WPnETP7NkiRoc8XlW/+Fga0KqdTPXbzt8XZuiK6lMMKrGcrf78qKSva0Je3Yv
FNguQNBRbjYiXo74pA++JozCMho842B69dP42Xn4VUNaxWrE1CmAQVtxL5yxGpZ8dEK5QZA7yOro
5WgPAezS2jn8g0ncmN8d03pz+Q1kk0Uh0BzS06az5bFT3CptIg75Hi3fn/JDaJbJZilpV0ckMe4S
aM/kkWjEoFHKjnuvOSyU7LIAXLfK9s0y+JtPN+suiUAyn2Vv2ZWsOpUSUDTqOq0uV1AMd2zzs7d6
BRnPkQqo6YAyPl1XKl9R/QZKJsDM8hqTTa4Go9PU5obCHMKQVpqR8fEuX8q0QjL0QpmKpG2C3bAG
vanMcfeb61KoJWVRPBUiWXoPlTE8fVN/+pMlM8uFVlAHNs3jsJJikxYl3GQ6RJhVIjutKqLZP3bB
RkR4ZZfcJM+Kzk+AFcRBB/3ipOKwoZH7yGPyt7+7kA9Xd7B7fZDUzrtjqCiRT7AK/rQgOz+jJylL
btrW+Kld7koP7hATMQoL7ob6SDt7/+yanADmNpMp+TFLafeFTzs7gJqmxqFBPlaVBXc/PyQkDNek
MfUPH8gAspuHCCf95CKF8fOV/6P+CopDUL67TxQRI+ISd1N9BtSJUuWiHeyN5epLqX4Fg1TFcWo8
XuJNe0rjtPkuax6Djs7d3Ive7WNxLnJ5G1ja7pYmVIKr7BtUw3i9bcYI2RbS1Et9m/5FJxz12ISo
Wc4adHvsN44/Ef4XuViFbscKpyNo8CxiqfNca9SWqxebQmyI2rgHgDTiIRpzUChU77X1lRSuOkGA
u0oAw03NwuvdEMhUr7QVwCLaCONTBrDwL+M+C7qz72wjKtKVSD3XaByQtAwZPCF6BxaTUIgnXaH4
DK8c50yTj3TfNPSQf7xOEHqTgsGTJMBg5br00DPW7UWGyjGbUKIxwzd7yUgNi5/PkpgeCZ4rkFfL
syUKlV9+1YP7ZabR0xDjCQr5Qw8SG8RBPIVANICyMdj1l1BKNsS1KT+HfY2wsThhwvSZmn0WLynl
l24GBuwWAhptNa3+vbfrikPWcRKVBmeDAMulQVs6BSVffX+y5cqfmA1uWjBZzAk4MP92L5p/7cDN
XpQSJe55dwPiLZijo6NbjGCyOPXMe3aGjqZG87v67T0EB/a74cTtZppwO8fR1WibS9JKV6HVAA+N
FoVy533XuqYchgEBzl9xHfSdAYuHcWciEojezTBqhTIsoQVFyFsN6DCTviurO6lUQfw3tWA0Yok7
C928OuwWX5baInN4h3OjVrVQ+r0xbFFMpDA+BtuR8+vjeLqeMA9WVGSdOYmT1YC4mI+eqZ6sgDhL
egNEaZ4UWHYk8i3+iJFClYHP7bTop3VmWGD00pZLUL/nTkp8udJHCw5SGEqk1jBCfS7oSLzVaNqs
UZ7zoiPnd3bv6CHQif7pHrSZbYNOgcF6MWDOhOtKVsPLkeKJuKMTN165VivUU9Qv4HxS9pVhw21n
mbgK4fzt2+LrPTTtv24LuSeSl6PEc5voRthnXatwOP55q+dYr1U6sBM3WB28D5s/FimKAAwE9UdZ
bI/cNrh6vRG33XgZ35xhxqn1Jf+mp+8JJ7/Vc53WCvvZ2WgsRj0HRqJS2VFHSgqkPkGrQ7wDCPe5
5Y75rHj3H6NrJGpkARLrshnVETty5pxXCDXQlmtjszLPazjpaCqa5mfM9/1TS7+yYLzZbnzcy3po
Fby7n+MyJCmiKjnCt7UNyRcMdKD4Ht4RXxMSFm/m4GFQJ7v5wRYQTftnUA0m70yZvgZhnk8VJLTt
jxajssBGcInA+us8b/7zwAdyAskO+bDE8XiyTRAM5pMcuAl4FFeR+OeWJ43xyidjJtmuoxgk9aRk
VcOcCiZ73pnvs+XISvYX3hxrY+lxFnbW+CGH2Kf83pDR3ZHNpCbqinrRCSLPcM8FqkOPHtcSFgc5
rDHnQFeJbgS+IiXKQXgdLnF3LL4fdFOn7opQVHjRg7PTRznGYy881W5BdtFIAKg8ATkOdaBWuNr7
93z8AbqPchTjDLY1T8dwGvMZWzIHnERSIhBdXhlfRPUpnW5YoO0XFojXBYxZaYTqgQl/kpztEwpl
gn5RvAjRuXCkSE8XotPlxArP3s8sxvr+pRxFXV/h0NU5GHAYcVVhOyBdx0P6w4c1tE0CtrhOBQf3
LdZU3ySBfiEHceN/YF+GCI9+UWo8uHWBxS4ZtYweEWB3qsvzW1i5cZgDtKC8o8n4tcqjf8YCvebE
BO9ZHZ4BZmjNT4J4ic52XokD+euvdcg1IxhkfLRVLggh3grrSC7+o9zRylxBLMvgBhcwXVOJZzGH
ug8QkLTQ2qnpWqYiBhF0XYaE5ozKfFXW2apXfxy8aQUVVOYAzpMrSddl/VLzN8SM56rFVnaURdST
mB+Pb8lRerDMi5AhG1WzatSfpH2XxSDp7ofJk46Nol/AANe330yc7BEC56gzR9N6uuvPTndCVOGI
WTpaTuC5vaOy51tqUXeFwZtEWzBgM9YtzS4wxRH+oxgOTVWlwAJ1B6PnHPH9AP2apG0mBWe9fKFq
I/+jy5fhKbea6KZez2kbvaHhLX5Rqv6Y+zz9gdGeLJGm/ZLbf7tj/GrCctTjYekkH2zbm25COZmO
Kms6IZynsGoHFHz3fmSMB7XMuK2NvPc/lfI6RDxvoCTaY0g0kB4ABtMtTUvJy2CUCY1T0W2muIox
w9/pIAzmaoU73nZcIflImVlCvi71byx2iN+l3WT5kdhCn3wpixddyB0s23U19mn+l4kCdily4y1r
dg2cyzo8VChz5yBIt/sw6XFYq51C8xMbdJEU0ZflBGpTJ6kFkr5masNp4fleMYAV+1xdyCUZo9XT
KrzqRbke2f9pexY00KWYrSIF0gDF8d6inoS62/OJQc43Oc8IVN6S0K4mLwZdFOVHcUGIwEg8QeEZ
1Xi5ueP//XdfPk1LRLoC8uhDykHpFVsalErBHruL8t/COw/DCIpN0f1rFaArWsU47lHyTE2Imxwq
DDFKcGoW5O7O6zDpBrsRC/1xRVwo0C9XeZbsCTlNUw3/wsDrOrKtjgHbbp9O5Qf5ygHOR/prNd4H
gsBhK7U1Z0SMaZstQeE9J9iZeoW5TEwgjdOeqVVM5lAG/eOZ506pjraXU8SG9/m2DHPVnR29hRel
0uUKXQKxiMnMK6hXAHGLVpJSXBMrrngSP8Y1CME7R6+HYsCnlqi1jZ9/mnbqhRyH7SiYVHOj8bRq
2YHP5zPJ5TJfAplMkbRCU1H82cqvS7cbxVU0WjpZHZNvEnoX1Jg/U8AZQLpQgU+xnhd+YJIxD4H9
ShqPeIJ/yWm0DriCaZx5OLpXsjAu6MEul2CnOCq5Xshdew5ww/1L56KXRBUfmOHJnxl6fwjliEjr
g4ythWuu4ekMzN8zeUVZL0TQ4imxLxdFJ3372gPM2O9gfwgzZRnQgmoOM4tsoy+6JJSPuTaH/IYl
I/jaXTxy8yzNfLjnpxcdiQOuQXbZse+JIx7fj6+qHw7cbZWXwFZP6NPMtbIjR4P5J9ZyTd1cbJi+
Bq80CQGoJe82OaEmOUnOQorKLkO+imt4fLOQCs3iYnNKHN46gpTXvQxyWB+44l1ROTDd7O7B+srh
EWy8fQ1FZqdIAeqKTkQSP2RlGP73mOqG4kr6I6AfcbT8u89+uTL9RO4ILuFmN+DTVr+s1U36oJ1q
3yDMyAwZfuojo4/RWkSlj94kRiO1whRlgnwTaFG02gbpaO/nkIXkeJgbusaMtgyHLE/Iru5CDWp0
hIoqyIL6hXeq3yOG1jD3LY8Tibk23FoOzS9m+mDdOorJEQzCFiND0Ffcb7PTHlsvVnCPXxJRtXtL
sxipjb26zmq0TSbcCDIAoWQqKB39l5L66blAtytkbCpTa3Tj5lXU/rbdReLikp4JSdak8hxeD2H8
uirY+dmjJ99Lz+YQHuqMsqelBnv7Qh4FHCXyBfgN183pM07gd9DKz0cEd/T1HvS8VNqn+TcEegSX
fDDaGfkIta+x5Z75vRtq2VvkaVfkwP6/Q+RSvPd4EvLIyWvrM4RHqYNLOSxDaMKYrFhCUfs6kmHt
ZCHfu9owDaiJeoaKQI7ZNCAXYR9DEWG/oBC8Ve/6vFPK7yZhs1JYTIiwtT9CwTZnY1O9Ep+EfNCr
QuG0nMW9CwoSRiERvi14/w7hh9E/tFADTCOTqA8OVT1wCxZJyiziVWnif6/IPzfBJjA4Sl5Fvmck
WOKzaJZKQSYbh0S01pI8F6DO8NG0HBD9CgbdWy/NT2IYhshxQr996h2j1bW3HKBhLYXl5yk4Rb4N
/7tXZt+scPFXDPXLnLfxjPZ57vhk8UjSSx29eZh3anD7PCsHcMFq3+NVf17VeV9LYkZ74ncEoiC9
jrwSXei+VlUtEKNKBU+ZeVeWjuvctBTHBVzPdgA4t7HhM8n0dHxecPTkuWzOXe1fbxGdcQCpipG0
LmhcqslcWsa7Xnsx6k1M1UMTCDgVCXiM8X2018kHV2UUzqDimJBQ52MWpRSJaqs2O6qTOkIJjZwB
K16YybCGcvLKk1lNd0ueftdjicowB3lTlIs15hYTs9kxGYNvbvOvjnk/9Sle7Me8tdABleezjDol
OjpcxX0N7hw7pQ9VCO93pvhMetgLUFJH7gDOrWyNLVV0cJymgSqwuDVDSLLvQjioFxRe+e2snxcF
UPgYzq0awjyOblBkhtkXEZ42S/i7O+GrEFdvscvxpgmBWG4qaGp7v1QZcnH1WeihwO5VdN2ci4x0
twNctdBUquDT9x44im5va0bWQmkeQlu7+vkcRcY6PTWuxRCeU5am9diI63VuIypIUVlcmDvsbEXH
iyH+ZcJICczOkiDzfYBTEUifygDMPFL/nJu5WoBr3oVk7q4xvJt7+tcSn6nsYQF4HM3+l682mNHu
qT5Jo/sCv3DUaQpn9WiL2uo9LbOdRj2W6JHUo6Ey60frSBibOPOxNmH3Vai9qjlEdinfMY56BzHf
qC7p3cyM59WTKRWuqa7zkF3eeGDFag/c23swxm1TqRLlHA5xH495h+GzHpF5uZiZweQoLyK8SIlS
6a9Whf4xOI+Vj7BoGb8c0vfg55RxHskPx9omedLDFAbPxzqyaitShf5NmXKummKUtJBxNlwyRP8N
Tu2aJL+5p4MqpjePLcfPDcQOD5FH1ErAa5jMWgjfPFTDlEIgP7RVeYON1LxmR9poyr0oofpOpOK2
AdG36JJ+YNntIilig8krgfGaV1iApPorMxjA3JE22D0tpztAnx5VDoPVUiGlvisFqHTXZKty43mj
RfEfJWCnapLY2l5S5G34YZwVdHnsaSirST9UHeZI2+xtBKFAMSmtckfls6Z7gx1SFzZK/J+xX+4v
KSdJ+8zUxMa2F3RzVuOWPak1sl8Fh1wyaQVmOTkMRcxpoo9mN6luJL9zIMXcNVzNHRmlpKljbXIu
5F2k6jMvTd9N/qyYWqGOwwD34tFOx3l2RtSN9f+UnVFnIXiy0GEuPJBQ99chjr8VdltogOwNfxeb
KCFHHf3kvAk6PLJ5FskijhBMj/fotJU+fQwZ/50sPuLa8tyHvfg6moNpNfijkYBfbG0C5AJgzvla
3Kq39o5nA2vk6ATVlJeYl1FRVn9T4VE1os+kxjcbe7D8PHWo7WZtEUSGLbvQGFpNhuWJgoG3q2Ye
PgILAbz30sagimJNCsn6FKot81NViWCJuMsz4KbTsD+35sSwTbMoMlPVcX+6AHAcRk+zUn85t/5A
JhDuhf5U8UUa9GuIpNUCwRsemUuGVOdvtzJVz85n/mdTgY7dNG3BYx3iNCslFhnMReIeytTIPqw9
n28rDYUNsc2hdKPaL+P/uUj4R/myPG7atrXq9oPTNMHY4g0iDe8l1Pc9+l8aByNiCZaYs8o6ZnPM
JSy5OM9KOY2oZnVPjI/xLV/hEPR3EcKHzwDTiNr8AkkKlzaLuMb6KIMUnJ7xqKr1iIJj21tCq92B
ZPsfkvB2hTcMG6TOpwo6VvprBbJsO8/WhsMYRpm6IcJC7F+ShifmRYd2w9rHO0Sejb1DBpG/DMaP
FyLaz1QmFSBYkjBXDyx1xTcnTqVzJQwVdCDT/uw9TCdDR3IBR9s4VGqlTafCHM7TafpDPfR2a1e3
w77sDxxKRcM/Vu5cmfi7f1Q+mkYDBNWQSHjERdc+/uRAGXpYkKYhRkrXvWlVkIEMoRsxgAuC4npF
Fsn/5kfMfjpsxrP1e09fbW5RTVFGrLNXsY+5PrZBh+rEJCHyvVb1SmOOMc6oCTmMigHM2aTdPxXZ
MNqpqVbNQ+4NmNinCWM8ZKU6hsQZyW9GtBHz3AkYRnaPyxTocnHrAXJ/d6ZOEphTkaDxdUXMygmB
b/dnT+XOkdyCvvq7sKu/I7UzLZiw0TmY1FasJb3kTut/kgXmOkSyv6bdtaJVZw/5KB7Wg4tXH9Mt
9KH5DbVYZizyEH2B2jWYCN8BhWsRHGVSql6Miy9qoUxdqrvMq04kauE0jbgOjgxmzljR9DWV0FT4
X3jVP2uFh+W/hD5loSC6ZeK8/PClR67s1jIpA9ofSw3jclJA7qwsrUWx5eUl9RcUI7Lmp12MViZG
PxzvweDibkKl1zeTAalfGzrTFfaC3/QTHaEch1CCRzrPvfCxu050O1aP5dfPyQBUfEyBA4oW4ERp
fXk/gF97gCbr2pLHxe9AHuZVXnFp75oeRyvlg2SVCyz1D8Ue/dBC8wHvLff4dvGXpQ1CghlYyKm8
AjyIgb+nJrK5OEU4q2uhPrp9eAhkjGrwmGVYvk3wV0NK/ZsojuxqZ4ivnNxroNBrgU4YJ6w9ig5R
RVnWrMSYe2SkZDudkkVbxP/oWHb8C86MApQtRd/kSfMXWuqAScxcfPt1z748YhjTJwfMk7lfXvTx
8azY3kBYKD3uqf4ZxWCHD5JG6kNDNstndorZQtSQOZssItQBmyiiZCPqcaEosJDKT13hwl09lK1G
1iASX0/LBnlbgCgVZWdDlaKnXPDGBA/NH0S8qJR12YmTaSY7wvjBKkMYGRJBfXR0QJhmKw2X3Vw4
bRPGP3sNWNImdFeJGYaj17XhQ6JsThNPgWQS1PLyc3eyUa75fNn4OOCzP7aWiFtDm2QLNhOmkB2T
qJcxX9oweVkMOth3lw/Kp2njlGzpULYLkxpJlNrZGZHP7ZjLCpPnb05XhKLh4lvXFhJfRIoaYfHr
ric6W5n7mOjwzalctv4P6/xBObBxccLebgtaVSqVu5aZ9AkJ/gSTWRSrnpBtk+HzTMgMf84uu2kp
7jIH0TEiod9GD/s+wfD6sOzEGQvZ16YvseniZC/tjkDczk94bPKiQwReW/+rizJyd5crjchA95Q7
ctl5Xfeeaz/RUbrXpVIbF/rRPpdEpFytd7msUePt5Vdgm/ItLbDw545fyi9/rAbkKzjbPs3fp+FP
3EIJ1K4AgqdSFnTpCT4JG5964q0co6pmyQR5J0xsP6Y+P9mQrcO3DR2uL/QPIQy+vnzCM/ZOLslN
FPtC7ePRt6R6nrPNuphJ/GGjQBkaDmqHudOh03n5sbWnWLjzCvxsy4/utraeqyLr0LJtdW1HO1tg
ZKrjlLK8C7Mf74dUAHsMgBM5POtkQ1oOmsa/1Uhl7Y//hugKl3/gSIjTF+D1mXr6p25mGgtcV3LS
Xe4OElAxe+3tlKHIAs9yVyoJ/IDT8LsYVkCx75PKbi64iifla76NIUqJwplVMF2m0vtXNIUNOq5O
frxSHaEPQMBGOKzVLmrvg50hzmcpOOav3uBp0md/xxQhJJfsN05CbWwA51UAhOy2H8ChZsub43ZF
DMJUbEY7jEdQGWK98SataT1ZYB18dl5pnyyHGv6RKVOU92ZD/oQXGDeyC1F/F62rQIXct2M9ovjr
WvnXQCHk/DuJDAlVLtVzChmKQR/tIIy8JEzh1AbYA6dWKOysJ6CLhH2RFN0smCqBEQRpMbFLhzd6
GOMjfKtqpgUwoV6LRYaw0E5sRVR7t6pKr0nQ02Y3hcepK/0gStU5Bnt6dPXRiMNOHkVGIkDNuciM
IukXW64+RGdyGVtOCNpBzr2nyIZ7c/YB048Oe2fVtSERaT+irP5gGmN41MSfcG7wFMkt7PhIFmDE
fXynvxrIQZ7/V+MMfXG/NA6145NafB+EpJ9+prCoGqiEN84m3EkttpsMhx1GAhqrNYAvV5OxHQMC
32/0KQ5HVZaDt07/Cukb2kNS8hGY4uglzKOzh5InDa032QLSdBcaCMey+Nkaom9JXyfT47EVKMXQ
nN89xk7M8t/9Izg1m5mzl1vGcAtrYzGP3hc54t8JqGZHOXRMCQiixllchVBa/UI0BqI9sqqTmM9a
/N+3U37tl/Jt0DTKDPehOJWsqB+1n+CVldvcIkY3UjAaBU6YOV7+fS1H8TWNSj/1Z4CVIrZIepN1
KL24IrSET1i0ejof50jJFhjSCT6N7FThj8xFymk3X5RoWw6iP+pZIh96/gFh46cjZbL+ezLAolOv
rb5DyO/k1n7WLuJrBtQcBgqkNkvpq1vh9d0CpZIppXfMOi6memaepr6fGGelJwGNAj+5KlkWydBI
pZOtvX17AX9m9LWdGu5D8vhmyb27MMf5vHiaErly7vNp0QJ1eHG3bBpZYo5z96X7zM850kCpp8tK
PP9zssJvN7cFisGrrm1jOYE/COzKqtTxtKGIbseQXGVUXcXhWBz2mosXS5ebMXqmfNGqmKGAzfUX
2heuKbiwEfKvdG0iboJhp/Uk8dVLt/k2BtkyoP09IxHqpQGS0tKjD+YX6lBM3Ddea6Xy7oeKA6+m
ViEuNWT/02lE2ask3HBgjTebQLBwetBXO1ae9yVcZZHJuDAYWbnAmeMwQT67ltbCEcIDnuCM8BnA
zw/alpzevGDhkExvtOXosxNoya/wRHssTKhthWm+Mqw0GB2GI3uHMhREo3lSOnq4GJpkvkZCis4p
r6Jkcf7qYpFXF+eXi8BUZVYd45XZA3zqweYMi/FXqhxUaiNZ5X1xdtVNiUnBRDTYQwg3IDVa/S9o
qHY4IeNweRuHHgAm68UOMmDXOaa10N4GXzE58KYpaE3+JI/OvbQ1+DJ0Bs/U8va8UL/xZiSEY1pv
btsjqabvqj3pPfEgKWZ9w6qxg1FlZNWy2rXnfFDmFxMYrzTPaQwWIUmSTkuKbRKa/FSgTKfD8xSQ
kM/2p+KFq8jYgG6m0uh+rwkSsL9tuGngS+Z9mv8UPS0fhUPdL6FMEIZSpS729GXKjrCZHYz0Poof
UErfI/pNp5u+rtwB5cZYSFgQvrmQnTH7EgGsB+xmX/uwk9qI4PEl4QMzT6f0ViRlzeINc/5Rf6lL
IAX6+0S4e/xMSZ4CTSoDe2Mp6jT1tNXys0dUQ2lnHhtp6+9SmLW6LCqQcnF3KInpIyGWwnJ6YeBB
cf4YGH5/vkm9g0BRoq1PGrUevSRr8XG63hSDDgZwByhKErowlkcYM0fZWtfxpClci8LgqhuuPwPn
DAbF/iQsNIFo5TRgBOToPhNTaYVqIzS4k2ReV5kZqOap/WP2tpnJTO8ync5a//lS33ooGzzKvjWY
Y827zzpy4FxKpPXI7xzqDEUyKql5EdU0xkaMCtazj8+aD6FLSD+Ak5J9guuvLSnsq6UIy5fc6Rxk
hTayyw40fYa6t0D4fz+BuXOMceeQTI/UM3YAJ299BQvN3iTHVdG477DMMwC58GcUN+1Afj37iVRN
Fm4/suCRI4oMMUH74Kv62Bp3S/xEwv21GC0CPODo+Pw5vi7+iqjVFwCXDD0cJoLqeWAxfSE1BhJR
EBYbhVpV7yzUxrkWiXXOHQQ1eq9IeXuYdlxGZrJ+gjvQpSmRmnrW20DnOBm6wypuaBt5Gk4nkjZQ
DmHhkGkpSvzdte2GOWgHjpG/grxfs6jdEx8J0VVe5ZK6SHheZRGbnCqZbjKFADwx+T0l1T7lr7Iy
JHvFR8EJPP4kxfxTz1PWdc9GxJki0lkxotNd1JibYowZs3j5+cXiw/aVbVc8Ivz+vPfvd89YMxs7
JOR4LmouVgbz8Pab1k0T/G19czgtHys7pdOVkCDMMFt5JwtEyQrGA4AdEe16XAyCRFhIJ+FplZy/
8ssuC1fVu1UTt4qP4E12hNoaJd+3e+O8A839vHx175j05FmRaCip5GYj9xRssM05+tf+JqL2d1iT
heY2Oo+2EMBIA+JvVix1kK/jwdbDZp1Pt95TicAPFFFwRyGHGBEI1NfYzeWeStor1WVq0ejdA6Lw
QH2FyId2nHJrb6rP8/DmA6EAru8ZxOci8/cfEPymGVo8CNny91A6bpDKBxwjTxZWIXMI6KbFlZGe
5gLDCfbBzDlyeGe7q1OKB7W/QuKNgmIx/D1jANuXBu9k4a55wCi4rETZAok7ENsHPFg7UT0mqVK9
yecVepxEU5y+hdu9+k0fsQc3y8DcZMsdib8GY4xWYIggSHgcornWTsaqJqIgpRXF8AdTN3asAjYf
S/qL4hDS/eOR9RnOUGKZxEtc9at6bhgCOca41PqCbyQYZjLPZcDW7/A51aNpdw4YMvrJGBl7xLpv
4iOnNjEgyEvOlOAvYvKG9MjKfOD7ZKinTy9WwgAgvLpZMdtMHvsLuPDVES42kiUCGbdEQNnlIriG
2y3hFmjX73SU4gWwl0ohsCUBjPEiYSeehQhOz0/3hkDLg8Of+pzIGnNxcSQwpFPoLqQJPiN91qb5
bwjOAzXgwPtT2wlDws5DrJ8YX20hG8gelSBNpOYfhKVNFH2zWaj2jOATwbEqrw8VDFWdSvashwEf
gdmOKzpjRf8u48R2BB7rtGjgbKynThE8np4Gzn034bKeIkcqXGk+KJCcgt28cQajrs5vGLz3I9Dm
hf0NCY7Ni+OIkS1zo0FAoQAslWN7Ji/S1kYkEnBjQ6i96nE5nOQq6EvlykMWmkwj3ssq5WhAzYtP
DZZ5e7lHLJaoNN/yUai6DB+90R3jijvAwuMiY12M1sYx5dUOw+4JF94AzcDgWkFo5dPDiQRGTr43
czlHajv7VwVxGnMdEYw5L/AZOHn2CMj5YzYnMhTUQsx1liTggqADAlNetB8OSjkOZf3IBfZbWlHW
rqRAL4lJEcYU//cMKlR/6hMpUznMmWQJTF8L4ZWFzeiruPmYHOrTJ9E0ANj5xaHRbs2mwRisf5m5
NlAYdRbDrQqCryQ6nNPf1KWcdgR2QmfbYvK0acIxdBuk1epFItQrolnRR3nN/+um2gKunsJ4q8MH
IIoNhoWKhqoUoBPLbjAynqu4t3eCPAyL0fb0ArRU6dF/N+uxCYD3msNYzJFWyozMYOhx1Tv906ai
bagreOzjuqgv2y3mCBrgBPvQge+S8EoQTDwnrW2VhVLi+RnVez9S9ZDdDZ4LjXbD5zOi4PEyyTmz
z7AOaGs6jgrQWKlpxnW8D30L44ew+nTHjKgtEdFfqQ3TQchRWaf+mmxIuhRrDDDRhCjGpG41fkXP
M8mx29PjE/5vipQ2aH6ZvJgMCqTtFqGrtSQTrszZSVwa1F7vv7teuh68/1DoCwAAB9VoKU7D5bb6
wnO0uYO44A1cTo5YSCId3NjYRMHYlmg9gxUTd84c9gQ4+HKuYz9EyptZGwi6HAmLtf6t533FPUWQ
CZz97qEiC6iS8Qk0zmUcWGXvarGjzsHRY+HKQfrO8vEAYlZY94jE4eUAEMn4fpfgIFVuZeC5PebR
uKgY/zyjbcaIlZJfo1uvkQX02QpXhNz0JSrJrB7y+khrqfEt1olNhnKzF+E+yYn7MDsKbY39SLZ3
bQd5qv/Z55G2U8uvo6a87xD6/VqpSTWnhUu+RB4HwK6+OSIFV+U01TE+pBIzrs6BpGb8x30qsZ//
n+UmxDMH6bcrCB2NplapBV/OyH0THszUr+zgE1ozoPMJAonz7IBSaoTezBpRXwUmcRoxDVG0+F6b
1n9rzxpVf1+iKaPxsjzzf7anO0LRGZz7il/tGUBkHWYo9SJazvQu/0CtwSFXK7BdW6SCBOIqEkcR
FwQGZJ5Xx/AReUlZWk9pUcyEiOrFkl1nYnDzs81PCSoIfyT7yNz3k9UxEwgqeroyyEOvEH8EeDp2
VVl1J4Sg/un6Hw46ylDbdaTA04sSkwOEG9ECJpWZrtdz1I0DsNyYw3hzE/cw6T23zqLv8tuTzQ09
tpZxPv0G1u3EC7h+Zy8UBfzhtmWvqKY6ZabUg4pU9CnC7MKwdFxQIXuPfUtqQhIZvcp+KqrVWnab
BhY+CtqdHhx9vWgJQwmx6YtE+HbrBumvNdJp8v0nuU883Y3toRhtJLmduZ4RxQwE58fqlyzdqQiM
xNjorARMEfYgOU7fCD4lpv4xMDnZChx1al90bB6vXr5qcLAonn8Rb2ZiWGZ9UfK7XKtIw50HZLKh
LV2BlaDysnQbs7UucFlKJg9b6ViZ8PAo0mIEQit/L6jOlVZNtQV49uCNOnibqy7hyBodzFryhlcB
a29o+o3hI+DMPLFvpJk7rDb1MJWej5eFlyND+dkDYgZKltAMT5cvaPLvIswbrbs96jnBY8kbOh8f
knywG9mDXUu98CPinPz9c6r4PXu7045UzaxfeOz+/LVjYL7oeYxid62jjxL+HzuxrY+fX5IsU8dE
OsaKaQ1TTwhyPCjwlCRsAg5sg4mAwRY4GAhdx8n9QR0r30Spe/25xX3hg9/gnesPawrf3HlhO5F+
hoT4eN5EK045oCCOuSudvVc9pQgdUN+OLWLlhOSjampU5cSviAtIDHFrU2XcevEnr7oTkH6evd51
s/59HBJBHfLDJCS2gX/Xyd86fCTAMSKVhyHM2tAH6m9WBs4Y9Q0prDMn29iZ8jf4SlsaWKGXJofx
l1JC9XMC7oKYHZQCs1C2QpLFfkK67oHOxo00GFjp0JLdaivYqgqdndSVAMafwJgjugughtm8vgf7
Of9VfvgB5VQ4J5M6gEPbXejjEB6P0eWbHc9eq6uKtvLj93Ou/447k8hzfSnEJnL8dzZ0rkHAe8SY
qmdDlobWgX5pO2ddtbv36JO2mklgZEXVEgAWbOdNMhLjY4elceFPphe725VvBzI09fbuukn5dTdr
d/+p5++kDzQyy3aV1QzjxPb4iuF6vir3csiF4L91SBwJ/k91zsTR9cALw3xa++u9qJKd0YPNVu0K
atchrH6VBibW2gbIbrBl/XNXnZ9QvOlnDiaY2ytUz9KkHHV6ZfjDhpYwP29v1uoPTWWbW/KgqcZm
0VeUj1BjYoqgJs2mm8t40ARy72SreJ3qy5QbIf+R2h8VbSf2cNyXPnnco4DdW4+qu/88cgzOb7Qu
WxVxDWePZqrbylAPO+fYnz2MDBE9l9y0IrHXdheYbd9htlHiKlp7IrACd8BVDh7idjBeMI/QqvrW
YEWlzO+Qla6L4RaGs3ZYZOcT7Irzuvc775+G/QlddoOczzP56dCsMJkiZDShTeNCb1Eo79tcs+bz
BoC4JcHz8AAtUxHn+tXHMwmY8aAC884Ao6Zad7U1DFNugt6r9zKTZdkn8PcuxX5xVAA+W75BY64i
/D5J6FCSBv2B7FSQ3RqY6auMXPBS/nkfQ/l1SfmJXdkSQvjQRfOKl62s9WRSpTrgDwOCLSrdR6wp
4JbApxSFeyuP7fqSI3jAVg7UVGRsLm2Q4LSEOuOiqG48kccJY71UGjlKrIWocuvlCVr0GN0UwHrE
ENYpCC4qNEaCog5bkiigLzNoC5GRUawjPAg7+xDdrye64qcO4YIJFkKRexcKVY5uXZqWwmlwBv7l
t6RMt7SiyNTycSgh7KMHq9dHX9jzfGRvcV5ngSZZn3nL2xxFPtrRT9YzzmwqHk9d2RDBsFVT7+EB
TWyCgfQRx7EQOxXGKCi68axtc8ufljz539YHa87O21TLda3MhYt3/ZHe/oH9nE4jwxI7K9qLtNK3
9KwDhB1Yz3Tlk5WkXZrSJ3XNFbruE02viMQCPPCmvLBUSpIzgAH09EcABFlP5FHWPRejeloe7TbO
jxYe2kjj6HEVcyl8gu9Z407s+kw6yYq57MB73+XeYi+bV/iD46V4rVL7Em6Gi8j0Hf826vi3yhQ5
F0U2UhMZ69JG0NUN5nEy7as6E/mETX91+Rk4fZSYLVw+ob+zxXtZhwSCFVKBY6E/S0WnsiyvTvkD
rjaNz/ysDO7HkHO17GikIWkCzIqZ+VHrkoRLSseJtfSo7CJpFP1dHp4Id63m0rx7BYX9ssSbDx7Z
4OPSH8nl5sIRlypb50UNT7N4xoNPKTZIsa4Z+HZbFAFqT3+j88xZNnuDVij9XKSwSSyfQt0iFrfy
jMpMZgVf6K/DXZ31ajk69METG4sXO8fUVCWJpHlcr2yEjoVk9iZrPEMXc6y7Un5wK57/iiyBHtF1
y0HQ06Ktj+zbnB+SQx+Xg5pxdzXzixwX+eBJbmVAvnuoiAtoQMtiSMEaI2qFZ/DVNPCr3vduQFgG
25D4DmPtRQ8MgjdyQDH70gsEceq7hnx9vzvAN+J0zMDhu7ZrOYVDf4J4f5w+hytXQ0ewK9aUhC64
MAUJ3UcTSZiboi4uRbyauL2PWtjc6PjhNLPVCCeBpmmqi8lKhmLMq4iCa3UuQo4ec1nO5/pkqgeD
BgEBgN0EqM6PmGzd8YdXvDsOAKu5LR+lnGtFqDbH+oA93fsHb2nfxFlalawEM+a7bEEBv69+8vXT
A7JpDyovUc0rpIyyYcBh/lyrYRTkJ5mAbuWIRsV4AFOyUbODx+Njwb62begZnR5307x+kEpU/Zfj
D0xQYZaIK6MiOevKMJoUFzh+TSkg1jxZ6WwN6F282NWpBYMoEbInKPReylxiglX02I24KRy5OZ61
ZwADbAhMN/e6ZF1et5pao8k9C+ps3+/2CVn/l7L9RnCApKrkXDyP3zYTak7yfFSVsrD4nTquOQJT
8HIzJ00aUqvI8SAJ/q6fBGXoTzKEP2Jb4lTuEJY0wb6dQum8KW3KZ62vFnzWgEGm8IuvYLjBosiy
NRJlbXFVjFQXarYbH6fSbs8cEH0GBELp25Rst0nLga26uOmlxZm8tc4H0jyuRoX8poo5MkRZdyfG
KV2/lHs3O27awFZGhIyEvi1KJNY+u6drGnmIFjS9s2Nmsxsziscb0QBzyBCqFA99WF3dzh56EpEH
fYOTs36LkGWTHm2JKZgre8U7BMsSuKis4lWMhgfDsWNkRODN7xlOuGJI56ZK/Kfh88FBOgAlwTc4
Tt/avqLftTiI1IfI/vWFWAerODjHZsbnRvOswk88QQcV0sUw4Tc13TulVgLbgsqOGajSWxdnSgKR
fMdexSGSqUAestaWm8qJ4FLIpkGlSWtpjzW3fjNxl9M6eCiNAG4Y6Q5HJNtHwZOZym3exrlmiNo7
rSVBW6ozZRsedpYo34NjWyWrK39xfbWUCge3I2GYORdR8UdHV5ZwXaEmdTztcaX9S+XUGf45Dirq
6kfx2X6FhYmoXjOtMnjrp7WS304EsCnjSsH9FQNbc6mYyNlj8TvySxj44dmFC9yhxiyYtrLSaVWx
PVcOUSAKEhWmwnI2kM9YwfzJ7VsgMKqg0GIno4AqFicDGoze8RF0TmSBPK23m+vLUB/S3YaKyB7S
By93+VDSTHt5KQwV3sPTklnwVsCIyse2WMvbhiXsllCwpajk1Ho3RWwOIfxdNQQZxFMn1YgyI5xV
IAaX5CLyZJ2e3PMJIEWYWX/JgpWYU0P67gJnRbGdg9NRmJIh1ZW+VtaqUoboAcN9vuN1/e9Uvzbs
p2ttcf/oqUa32W+IywK89iIj9AlEFfpd4YntsU0AIrTWvbA24l4EuuR2PB/waeYQKlL7uZa8zoDy
1E0ltf99Kq6/YRdUPAdhd6N4QNmCii3b+yNXmqdzoysjzyVY4pOZdqpwuonTTtkt8TZ6iQC+7KwA
ASb8qRgmStMCxvaQ6o+edu5RgvtOOR1eYsRoY3B/WopWi9JCaeMEaEtIc+U9FtI2PreBo189gGny
k2qfpprAapxT8168chcK5YCiCwKchqiAwWnRZ76LJaMLNZg99vzmxdfLAvy9jTITP7I48YNHW0s2
Ghdad2/J4H5wUH8l3tuJWFOA6ZqTkVPAl9dBg0LO8Z5cimdiHKx0km+J90wSJPFvDr+m/rfgLT7e
jxAyT+Ku7eauM5gGbN9k8NVdgFGtLo2lqLRdqCwbPsrsDN/P+xM76wRP6ciHWKNS6tM+jmqOsr9P
W17P2MlOUynrpgHsvzjm6uXKHOTgQq9vysDfQJOJyPrrXGhIWlx99wb3vtxFpzM43Ny4Tq2u3iO0
Djv9v+q75P4jBrErehoLTUVelZ5CNEWUyCG1DnBqIZnGqaJ1vJf+igP8plVwfLXm2qeK8NGns4Gc
OS74bB4A/vUP3EZnbzs1zTo8G92kXzLrUiMCVdHsDy8GYgSvtNN+XnjtNI53EeHSdIGdWlqCL+eM
wohDahTma6SE+2qbZno+OZiRalBDo6NqW2emsph8D/+WWj5JJ4VoWd/c5mLBKm8n8UJ0qkNSiR04
0BpMKRS7IWVHHH9gN8OyBJkGFprtKp/isxewQiRMMxXfsXGikpDOpnM00H26JNaYWu1HI8q8lk6u
tsaW/+CH7cI0wkPEFlR68kwzcBQC+6l9Lw5+yB6C+uKC9HgvmAh193Q8ABmGKOiZL2xKAmsx3aKb
2wP8BNyZ8tpQBKfkf3PArM7o5IN+D2yHLZQNaftiq1NWvyb4Y1Sld2nUJhjl5XJZqwpn5B2sN2x8
WHn6h0WDOOR7ZdsVgeM7H/p3HkeaTmN8Qf8qcp/Eoc8+lEV/8Wm2FitdMwXXPGbWNsbRAPyUvP7o
BOmQhFioO0g7dUdeVbugUn/KvLMt93eqngvhWhsp+PoxBqNgd8pE7Dw8JsI3T3Rk6PVAe52OEiCb
fuYFZg6ZBJHzCxjigRye0QXLfmIPW6XOpWnmsC1QjZBafPKuqHFt2S4nACGmRy4Z563IZARuQN+K
mHnxEzYSh5nX0AKvE/QKP5HuUCBcuuoXIs4/fOWBwBBQplKsCcDKODVhFlZzQzM2OBjLk5dOQjHB
NfOoFQ/mmaNYMMPQbFCZMtZX8v1Vv/law+bU172GTUIEagiyRFvLlrc0ZYWfXOhj/6xKMuzrsl/n
pEzZ7/w5tYs+h4OfeUQieFSzPVcJ8gJDTZKdU2awM2WviKBk1C2e98YwvJbNZG5U1Bho6n7dDL5q
BYHIMD+8g8UZPzEO9HS0m8z6mFYzfgD4ds29G7Dt8NAGnrHPIng5kLCLpUmBzTn9Da7ZjfWo6NMZ
eXwQYtiUARm2kTDBuMEYAQaQckNC24XHiarpF3x7Yvp8UIi9YKPl426BSaz6SMgiVQ/nP0GGiqSN
Iy2QUFCMmtp4kiVeINDy5T2mbuzKVJv74sTxB9+XOxJop7KgGYp2GI1/4/RMhehvuQ53Ch3UNsp1
by92onTX2eEtM6DIlYJ215A/fCleqdIWThSiRucz8yUyAxTa2MvLFhPDuEFI8oLk8QYuAt2p9tx8
4qjpiFX9YoqOnraU8mSPa3LvwWGuv6DYw4tHDX3K2dwgLqKSNGoA1/ckvLyIq7vuH82jwtX4JFrs
chD4X/vN1wTgwbJj0S2VFNtkFtAMvfeKtomoVMAKic1Sc67tnmwOQYBg8Z2M7VuyEkwgEbAtZdUY
ApR1FK+04Jw4XFZEpYv1kSCMkeVs6iCX3UIeIuGjkWa+SL0+gDWY3Jtz3KaTdSYytqf+Row4twOh
FIn27EYYfRbEd5aV9NzWTEtco8/28zDGQH748ginXbMi/RxCZgi2EuxtxU921vQ+VBSw3xsctJxS
308C1qq0w0HYdZvNpAcP35EshBG8x8L66isoRFVXWt5Q9G2szORUJYyYEhQVcpg9TD/Uf68e+CQx
8FNhbdJ1WECsFKG9SlN+5unmKQpbGhSqc/fuNO41Mw0yv4byRMiuLJnPMFq49xtpUkqmhC87nPie
NMeY8tco6zVpQJfUc1xNIsSDP4ElxqUNXI1Ik20muXQqZmsq0aavQPymGDNi5xm/Riqi701rghyM
Bhw1cmlm0kq3t2/8Uwp3W8b6zFPvzkT3ojJHPWSR8L0iIN86gLWfuTOgCOm/8GgoWSpXhrqVIXYk
zuaYe9bB76hFXUWWKPcpPbJbGrK21YMYR4joS5utaZ9FVVA3tD4NrlsIONzmemhUQ5mSeQfqdaCq
kVcOo4qb3nr978X5vCVFlnDc3emimV1ut0ymEJX/XgBi6ECdlG/AScMF1yTukoOUCEbkGxckZoMm
ECKwlynD/HcP/rg3u9AOnZKyk+ZOK2TEOH06q3TyJCONC47O9PX/JqsfSpuAIEp92Ts0wq9jCz8T
E3l2bzhFJzkvyzgJ87JyNN5Bz7VEJOln5XLHcrxw3Nr6SjfIIunUWvmWmy4smrbaG9IQ/3S2v1xy
46ucqWxCx/dAAKBoXs3mK5dklCirpH8bM5M8WOn0ovL+Trt0Z9h6aBslsqybqxrjDJQJmkC+6P3s
me2Rde7ZmuI+St5iADzpVExihrEypOOGhc0MlwGhYrEHA+xjFJ4sJZeYD6mDbp5up6D18AcbZfTj
s7p7rhQzTmXWcHGy5UfJ2y+q3jjFHRTnhop7PfOGd6vK4WuktW1gk9SV9KSHPBnngdNyDOFhatJB
npZgVoy3eo4lzjdpI8i6M06KY/w0xfdVHmaAKOVVKGrwfMfXBl0slRVcY0BZgL9U6Wk/FU0Dzdxs
aO/Z8GA0CEU/750xF/EHN9TFXyFYh0HgnBSFa1A7se/+ZUyKli7s6DToLHrf14bYgpitoQH3VmdZ
o6/5aKVfRXfI2IJnSStShRqDhLygTHHJosLAylpkMJiOhkMiXBtlR+tsUBO73Ez3HnqPJPIDBYmY
V6LgTd3x7iACFhjxQUyVt9CnyGVxGTMl65Ac++JF+OgXC3aVa0am4vSuk92XH5GBGIiVJnMMPqeG
wTRgUwbNe4HN2ibJqEqOBJKWU50Vp9ayK/y5yFwkcnOahnV7bj1Z9b4X2n1LlttNtDiN20nO4H0K
Nuz4r4+Uzp0+iCQiDsFUWl/7x93TPB5kqUasG+Rj9YHSYyPl26AiW+n2Vvn/wwXLpmZWwVyx/iUQ
6qoB2ZGkh7jMcR1CJ8nDT6YwMhxyKOwl/LSHn83SVE9vqoXbugxrV71incaxpoZZpB6EpMO1tBe+
LuJV2sUHEwg+1Y4sRAKoczC2pUj2YC8gy/klRlZOA8V+0GmM3BmXvjC3X23dgv+X7Qbr9PYvKKJ2
/E3E7pDOhkpxH3Xyrx/ldI5HGAYnzcsRwNMzbkt5hUmRk+NfFGY0kiNhK8Hid9vafHEJM0nH/0Sl
xRbTkOnRhL8CRzYEDNIXgwvqe4rlyPM1H14UqeZUpY9OG2VGsG8EFkn8eLmz/y86TfPIn4OEl8MQ
596CV16/lq7rirhEVqXMmxoFKuZrr6g0LAKC4xSv0YTlOZTaS0rCLGvQFV23TOrHisWATP3mp30u
cuSQ4ZQUqUrsi1etV8iV4O2LYh2a/7gyks/hc7lL+DywpSYTw0/ss7oR1VM4igH4AOjly36Fn9aj
q1ByUZVprs8AhnX08/00dijDC18KGxX/xzulA4ZfggwRZIkRHHjT3tr8zzL3FTQ+l9RPUGsuiMOZ
bwgQIr5m7U5OnL/oZEx1HaNmmoDQpM7JZCz1VUu4PDsblQWTM8EThQwQLZKEYWENwtTm6BtHuQiT
DwrUqYXzZAnzMrOav3b/QqAiu9NB0domVzBXR0Te5/uDm35AnckGKgSjJbuaUq4gg9OJM/N3NFkh
CkAQi0WIpZdgsjGcZlpiDSOGNdQE2fPkej2085g4QhJIm3jLYF1au1hmLVF8J+D9LnV1NkmakzFK
yRos/+aT/vcr16Tq/3E6cumgokq+NjWilUqa0SUeyYLlnh4xgTpEmpkzHA1/MLkjOLOeirJb/njt
z6O78P+rGSoO+yWnWHbRpOOvjyMZMMg8e+aM5mBfWTDKg0H5Ze828BZ+awkECBTioKIPUYuwyr9Z
mIOdtEQDhpakuybsZN+iQGaxhk7xZJDyMpepj0oNBIJyyl+HReabR8rgwHW18YM9Oop8UjSTtvpZ
qfi7wwONhrhggyF7qvVUSfz8lj50mSDsuHc79bvnQi+LZr2acUufGqchdkqMVQhk/rTk2pvMCudN
JHNga8M7iVDNUiEx9swdcopeqPP27kzlY1WJyb/3v4SpmEm+GUxf+C+orM8XbVJPDgUy8WtObHcf
auZR99ausk4+1P/1hm8P2LbqhKws5CHYco7Lv2jDBP7t+z/Dqa32ekmIVLVAxWsaUQopr1sPlrzS
l0nX/kneoo0TL6X0cZA6vGw6rRJBLGS5IRmW4+drQ7gx4/iZJ+WOWYXKVSdEX8RGVMUxhJ2Z5j0c
LYkJLxD4vva1VBbJFdXaHtB5qKE8BnT/9AQoVkjF0cRvXOZppZz6Dtk2XzdqP7MJQOPyBne1stFf
HEFJ00TejI6gs0+KLADu7OAKznh9BMLUzanGbkTNiEvd/WFhVLOzdzz2l08reNWvwEi2BM27tBI2
i+EMKb6VwReag5qbz8I1weMlZWNkjBvCPnCIDjexYqB62j1gLOCk47oy8VfUA3N11zKGqdRCTrkM
t4obCuLGDHAmdbcU1MFhzYpSHE55n+MMKHHHjQLZEzK28F9fPhGAsmxuQna5vzPhLefwsunGrrDu
tJSSEaqAUcmRm3cwNW7izWZuyD9QHXi0tWGPP71pI/ovw/qimr7KAjwujIQ4CsBO7iPn/aA7x7us
K30zLsDfTFN70xC4pLc/fdkbOG2Klkma7ElTNsJHVS3S+Vr0ezrGX1McsQEGcTZ1lzYBVtvFExph
UHXOOIcubZYrTVyFdEQ4wcZdw3hk+sO4AyTuJs4I9esrzZ8Fpo2hvqTr4oaN51NoQqPIQJiP3Ylb
q79sWfxS3jk6h/Z6Lmm+nV1KvSMnZiaDg/ma9gDGvDGtu4w/S7FC60BBnLKI3qyZyE1DbwlH4bI3
aJIzNescnuKw8xECgdyYRIiTHu2wivKRU4l13kZKRonqAHDOVBs9W5ltb9mMkVdtGPz8Z9lSWJIa
ESsfubLEOLvzlznMu5JE2VHk+nCFX+gFbbKlvVN0Ab70r75D6Mk0IcKVH9+S8/Jov2TJBJ8AJOZV
d9LENHi7thMVO2XRb3QARNLcO3CR8YlUwHFK8stLKZqo43wGAPTpGtj5NIyusrvG1M5fiD9ctjZf
rxXh7zx5lM97gE91YvkFCyhoLZNsWLOk5cfqdmrmmjVevQOPydzP4d6F498+IHi7YdrrCcr5jZSD
ZxayOly65e8i3JoE3joJ4dPWAqUXTA7ac7NEJ3ObZGDBzudp/YtapXeHKuxFoCe/v8uhseXRdE7G
W7fcR8cYaA/FZElI4Cv86pl0PQRcSMtRw8HWQb0fUHeBpP96JCse+CahdkcxH5SGjFrJVi+y2zly
FjXuvzj0NYdjMZBlva1dVWQ+jZJVxQ9+wRlohqpR/IlkMgqXIPf19P8Mk2ngZaEok5Tauy09NZXN
r5L0I8tRbs9HZY7F4mYgHeWjPxiGVh1U8Ubv5lGcc0k9pVs9qvge9xWTmPwh+H7ZI1G9CO5eyZtj
sJDk4MKPj6J6hV+MSC5ZmC3Ct9HFyGM7VoEFzCWe8zVKoCxwWOzVPsZO+MiS4RYHHLBPqUQwkqeD
JNKfC+3BVMbCZT3gEVpy1i6l9lH7i1oCVO2FnmEO7FSXQn4cvTsjaH5HWRdIconwypR3zDljmcFo
N0WUrCYH3pB9pYXexfEaR9DBazYNMlszznjpDrRhV/G+My2Wv1Y9rJO0cKdKjm5+gD26cpZAGvXS
Geq26Z4tSfOFDgcP+BSvmSsZtlwFpO7PrwXnmBs6Nc1Gw2Vaf7hppkj7Mfo/nS5Pjghp2wnwh+9r
5jeKlsJMttHV/0d/33y13/070nFrt09AdsbyiOnNHMkxHZfWnZDWs3A/BgQMAd+OpM5S4bgZigJD
ucAla7hCntlDEyC1zFExjeiJKf0Vg7P5h16DtBOZ0ChAupdgR5g0kVTldsmgrA19Ub2+hx90oUER
I+w9xupjSAzkYsML5PslQenEo8dzZkW4eVV4QqBTzwDVShVOxnVHPVRML6HKC2nHtHpp+G8Yx1q9
bKx6QAKtZIwrSaB8feOGv3l1Dt0t0Dyz/jKARgbsYgjNh6ghZO5qVXSkfcX6gojp6F98R0JHsmkJ
7h8v7Wk8yFKyCmikdYo5Z9ObQRjD1bepd5ojKmbKQqVy/6ktvp0umA0ufka+cv6DfBhTmji9zWgC
M/k7urbXPjkaIT199qLhRXlFIEfw1NucbZNYq+DMW7lATDEr7V+G5phYMC+FjvN2k6FVJcHdybHi
SG9QiK8oUQAKXrbNrzvOtQb466GJwT9zWBgASAY6vW56DSm8YjKGSY1t7+fbNjOOy+SZ35mZGqx3
YviDbksL18GxDYTpNAenPYArWCgAeiZ/dGa+bYUfSlgnTt5StTOTwQcx3hBWi8CDqBvYoE/uqq/S
r5kXehfrqp4BVqcEpR5qu3zQpRsCmXf6Dm1vr9gltuM5B+l9C4vuTO22SC1EHwSVJTwxczm/bZSE
gSvvu2CYArWunqXZBtZvZKsBEy65H0Wa/Um4x/yE3peogUG7V9Ped5WQ0fG2zHghpMcdycrs6O1i
380LwBgbRgU5ACDUtPpz0PIZOzNayAfmgLUIqYMG+PtBNNECErA63X0wj01KCdiAjhl0v3/E4/k2
557IOx2OoS0NDL6eSeLhL0EX2KtPFo4FQpalGcL4UAe/mVb1pZZfjwDf6jJPbPn1wswjEeej7G/X
NK4649wyGHiKsPBH+jkdFW3Oqznjk8vujrIT8zBbBn9+mjBNc/EdIo4ZZFawQ0WCaTvIRsws4TTu
/F8gS2UirU2L5PXSEIlwXbOlY/4xN0sPlcklvWcbQCloA1kyUpJTnabawHt8+aG/bxp2BqZx3raz
7x6He01UfDtoXLSLDUjk86q900o6/tV/a7o6bVpcElFzgBPds9mXMi5SDsk7oJLgJmY7W22xnPir
RKtRkit4b+JxTWz+uhC4j0JIqS0y2vx2ACXZUkU7q2JdYhij68kT0gcxD+wL+So9wjEKgDg7RzD4
xl8SoD4g7hixU2tBnfnC4/NrKA819YYmz9k8DKjs4mtgmcJ2ufbSyM2OzJ8yzWeu1iXG+ZtPaJg/
+kQNbSXmI3OzUsUyfyT2A0j+t5SMgW7ZYP+HMlKgaKdz0ZXQpWG48h6NPgXYg4/tu57Z5jQ82CdM
kvU7QjCsKqU98w6XVqeVLVM3M7kNKOKFeI+O3pOpNg+qzwKRYojeRccOxvG/d1NQis6/QUTw4MkR
cBqi02uyq3/wSR8ZDKpxLSERcqD+6Ye29/OvuQxVhyp6C4YJ5msJ0e5FTX2IenLDgkxTW5SFQijz
Y9os1nmaMdl9TTgYrFHKhvlmnObUuGpE1bICAUMaanCIFDbRG6sSvzIQO3LBrdqYauBmnExWqDpW
YXgrT9WeDovyAqTLEN3rYOzZBg3OZL6UVuvRATotw6KuiUrV559cj/YtUokFPZDpB5e1dEj7N+st
UMA2UU36rRHnr821CAmDUxUVSkzt5+aFjaU6KEYgQiOPiVSusQtmuDQjo8iv2RzdFDgijrMpYfdn
N4k0NIgQ1iO8doVpVMCzjfdGFvYOWC/eY1NUAfyoz9GH6QZdrb24ig3XT0gTyALgCMpTCjVuaIuF
tPZ5VTk9crzk2dD6oAX18UUp2oiPY8hrMSIVlqrxl6e8726siOluSR2XXiil7IjX/JbiDaWlsMGV
vfN2gcP03gRXNuw1ZQ5D18u9OZsGqwnPtrV+gxVHQn4tCXKUrH3GBc6wfdJMG53DdXd4WtN/jbPY
EPAellaQp7Ch3H8oWcp19IH6Z6FBA8nxD/OY1A55eGMl58KSM6CJclHpBZX0dO4tUQHNlq5CM8v5
I2s20H9+Y7yJ14+fjpSZfl4Xba4EDVDfaObm6zNlSdefhPQMkabaHQA2P4BWZ8EPusxdE8HDrIvR
VYEIm+iiebDzpGg7lel7DrBHgacuzzMlFyKUcRx760LNZXP6Gr4w4Pcm+L5EZEMI2gqNi6O/LgAE
K8d5r03xOwKvM7fsyjavACFmtD1Qd8Aof85BO7SbFStXMU0LPgXWSsyjnGP6sqUYnms82jQRcJDd
x2ZBodEcjv8yt6dGnOckfbvGELRb4Id/pnFc2D5BKSilgP8/F9BqpSi0L5L+3T2hBlwTF7z8fQy+
JecraOT2KOV2eOBVYu427K5NsO+13xov/9pwkynhRr2FqTKiThnrZFofRZg9En3htAit6Db5okUY
zCh7bZNER4GlhG2ZPqNLjaBjg130FtSIJZW1C7BBMdx3aIGts1tLhPVtM7ycnPf0YqmQSQCJvRy2
QeUzRmkfp5AEef5uSoBfRbex+SpUaeZsSpxObcFZoE/PMf1NhrtzXmCUGQbMmTDXCqroyqfX4l0i
K8t+qXOvu2F+2HSM5PTRSJDdei8OQDTC1WyLU6QyiERENwdQV2QxMZRoxabYIvdc/o+Ubx7bc/uO
yyWzJrPCY1xtfhFiOQsxE5AJc95EP9kKj0Z1aEk3s74J/4vSM6ey6Cz0AoDqWn0RerpLlw+mRtb6
Moee+Nxog0j0/RFHPLyQ9gq9QZwCeZ7o2yKlNJ3cqi5xwhGrYK+mvved7JWntLS8MFiJjJjwDYlv
eVQfot2brKuEcJdnkDUH/uV1DpKLStoi0KJcZrj9p0nuNqgcA1MbgBagY/Y0PxFMEy2D73Ny6TEX
tynF8BPTP5ArNuH2O11LpVrl7aBiV6qG+FsuvGV2gRNWxFMmZlqXlP4g6BQ+kmSDA9BOCtZ04vus
zdzNCFBGWbdkOwvSN5L5UixAdH1J8PKpyiXKrF+Ehpy+5Bg8EDTChKPH1RJ+0zcGTNscdQliLuYr
oZpf0DHn3Re7wbaKM7hkTilJ/qP7K9QPJtYR9sVnWMEbkI0gx15w98TeuonYs36/3MeRoMMPabK1
2UMlU1eclDywjaJbIpYRkoNN0oS102i23MGiSf1DgdpSmgZWIJ+r6naF2862XKO7WyXHGmTltv+j
M884++bJpxhUh2SDfx5gJszmvaUDlg5Dae6KnHAlQ0352cpWWTQMKmojUVZ+wGCHpyRsPpVTCLIX
ioUw/NicUX8ZPa/JlLJTZtla4EIFxaNDTsf2Uff9WI+Lu/qLFRy+2RWiRYOXmNwDjs/4voyYzpIw
e+fDE3iFn+iPZOyDi0y5y2GGNbBZD1niaVNFFQadMUG5AXQHBiOD0bYBen1s5soHsnYWjSkO3Zf3
DhQlXIdBHUBRBTPYIAYUcTmjzcYvvKuO91vacUuEeaI/TScU96j7bD1vuLEocN6pplmOmb1CoKVb
wXBjXxe+jiB3Z2H2z/oJUzjp514HIzobgiFjlbX4mWJ0xrY90JAKIXyP2IpkCkBKh9UxYIKMSIhe
AoBF55Kl8BV3e3y1uxw/B2NXzhvKsrDfoJ8AgOcHqjDLu8Oj+2TVkswxePgA5fuNviBrz32WncEc
jNQkACSpNqUVenIAfgAqdn+YYuq5jIWpGYKefdg0M6MMDCRoKNIv3ghMZKHKae6zA7gJq3wOO456
AmhzMcLN1j3Zmc3qut3423mcLvcqQDFSsGRsK9SY/TZXgyKKhtlWsuhVOGvg9Bqt7gwtTYRLf2ZS
a51occwYC3jUUmRrjdawTFCZt4GNA4kTAm0HrswRDU6R1WQl9avBy7byov/QSTEm+pL2Yox5+YCc
Hg2VFAvoFkp7gEBF+7nnCMzDm0DCjjvjH8v7vYAJk7vPIjvuofCfzMDWnUgtJ9Y7ooQGbEOR8S6L
zFC9wWAUTp3G61aCyz4663b+Q8t9yW+Q1e29J6WeurlNrdlHJJduv7u4fslGQg85JNo2hj2VfslV
pM98Ozc/kpKyb316KhwRHWvzleLYesS4Tdp1dEpg5hhlD0d8eHeeD6CHuo7z0GJ2fj6BQVjiuS6r
oWEt7fr9JR3/LWe2fD8Iex5EgebyEZZsuV4MywNfKVEdZlN+tinZFwMMwJL4Q6rCVWGIuI8KF9p9
nWufHdepHxtUSJ0FHCapbip1Fd1gFqf4s9wHly1wAR9JjWZQMSiX60h4B/N9G+H1O+ZJHzNRhQWe
GFPJDc2K/yec42hCpxYOccvlz/IJ3f3eAT3IvEvu3+UM8oviQn9RvnP+33it0TlFbfbhFSE0byOb
8vqTDcEvXqLtVARNDbqgN+xZlalVWJpIF/xBhwHRL3ciw5la2ZFNswrMB/1akmaQPZJ/2yUzIHLb
gnf0vIpAckE+PlnaVo5o+zbEDMewpEp1q9HmZGT/KfYfWS7OGwdZ2UHllGJEV2BNSnNp6FbdsmCM
8Hu8ymf5UT3jmcKnVwQd+LwUsdAKYfiSP27YbzRpk+xtG2Bw6CTZoU9KydHMEqAS7j581nZwaXSS
Lcf9BK4lnyZdsj09oc2wF4ZeNo8O/y4XYk6D+BTsuzj0uOxfqFtXVfSuou7ifT6Jfae+tYMTASL3
PqrPfxwL9mE2aVLThXWtgmLor97hfvLUhPtwr9OwVU6YxIMfCXNx3MWQtRS5S1b+TOuLcVZg1fUD
gRB1HJ+7ulXzq2YEdxCFXjhpH0rEaP+vlevH2MRnnrwagE2Phd6toUajsv4iDRm3GPVTYmhxmljS
WC6e31qJZLWcH+gq+FcbW0+htkG/5Yl2eqcflRaC3O2qKG3uxTZ8gh0OdMpnyU7/cRr0izY3VtqM
xfO7GmsFURiTxG5Yur0FkEDAv1GrsWRL7Fc+/gHh9yUzZaC1sT1Oh53bEh9qbAi+CAUqlKLMjn8g
m8OOS+LUd67O0Ju6wBmtCknYXlPE/z5ha1UvZG5k/0oAt614ouUx0VBLMXA7QN+5JgCxFoKgrWN1
6OLkkbX+VXLQCn8dM3lRcFvaofwv64q5Jumf7tbpYO5yfFD7zD1f0TGpv8+qgSwdAZJXF2Ppy2WS
8ZabXX1jAHsYvf5TXA8GdoUSuRJhk0mnWKRDqQcT87nNk1duEEgVe8iiclwxrirTn86CfXyWNS+B
Bv1ZDQprohWyaqGJTn8SivkzIbah6/DkZZPaBZHccGi12p3TiH1/XjFPJrpJhu7v552zot3fyAPZ
vKcO9Lvh1ReLmDyvQdcDOapPx4+VA6gCC4rXS7wGABA37V3r7nOM0f0ki1BqXYNboG2fGN80oB7V
8NHg59PdwMlHcqfGqY8n5U/yu4t4GZcFbZ30uGrEoiWC8nySQyrZgkzkfvUdDGyuoKL7bLcn3wYY
3XwN2rFXAnU7EX9VyXVR3k4r8DjUGL85ZQnjETO01/uJk1nDUKacHRMato8fi3hcl3Txqno7y9Q0
3EHm57eGPPOyrK8oeqDzVms/lSmqAakyZPMZ9E7ZeuvfV4h7yUhW1HdqrM/D/qqoi6/eicFE/3Xp
dlxsCx1/UK3c1XU/xrAirFLNL1vMDyuEeGShCpPs2P40jTuwwJd2Fs3uUSilRAO5xbLyVWcR60JK
1/9D5PlturKtqL7q/crpxXveHcmIgPuXL/e45jYQMQkiP3llQupPzp/Lf5xgbj9UE4rGgamp3ZzY
2WONGAxD94k6fFFkfz6LoBbE3U92Qaq+1uvw+vZMBKsLRXt07LE1xDrFmXgX4VaxEftg62EGnqXV
YXWVcGEaOLAivLeCn1ulCEF+yKEhEf22UZXcTiES1iuV1UYKc8e3dmPnFEms+ngS5G8HfgueyVF3
c1SJL1K7Kf5UwLOoEMS+iw0u5PqbZB67wduTgIWWdQPHxd1vyrbhGN6LGs/oEolJW7rvWi9zTrJw
3yMiui210F7bPATjUqpRjid0KIsUI+2ZEj47EOeP4nyf0N4z3NddCAU9wiJbGV864hOnqV+TTMAc
Obb7IhdEhUueQTHpsKfgiduF84exnimiq90baqG2CYUYREpcquixA8X3ehw/ThqG31Ohd4PogM5I
JzHYUDnFtktyKW/W2WgA5TlB1Kbt4H6silaXWa/fR0wwgrJTyGLYCfDz1pQ7TyWWN20pO7ZCPt9C
YWBAKLt+IoY6TUE3xezt8w+2iwyq8EsnMotJon+h2cnuJaYbUWLoco5YMqSJGd4OqekSkJtsugmC
y/LfqzarzZFgSXHj1KdTsyzHYuffkYNyCU3YNjZsdc9E0xMQkAa1w0rSP/WKkjVE8hBeYfuRyjuv
OGPJuXlubZdBz6odmxkcpQAC3QDU3jwoL52pvNXsJ5UwSZSE3+Dwazfy0s5Uv7Y2NUyE/b0vOAUS
3ibgTn4ZVYs+EV8g3+rp76akYZTSHjqI8gzJ1bgWKm+POjT/LPkgOu9/DMfbH9ghnN7hCmi/Qh5A
Ixe8+BnmpDVvzfewfPol9FvPwKccrHkUSwYeVJ35+IWpP6yHyiOb20OZV+3u0N/lwcMHs4tEj1Cy
ob17A3muoz19mMV6IfDE7T2dQdsZIBybDGLoZOXJ4MxayQLzBSthPwpFQN9uh2PRU2jT6tV52FP0
GvBb0CnjznoaxB2zJzFA6tG3YCLNtuFNEU/lk0jBcriQiZslwV0XQxmTVxernCSarwvyTYKSzEw4
cceD6q+GMQUaaBylzg+/RS1a3ocIifEEW34bSobsZo75XNPXdLQLPpARy5KVqIEJVb6JqHBwP0bS
MIj0OaLO6cwEbepkK9jJpcynLf3qTpN7dsw7ANRdXIrTvPq6XDzDFTv2NqQ8ocJD7eaucftic93n
MWxP2KXn3Y1aYWy66lpdDaDWp+lsuw5HVoMPwqmO3B6y3lEZJDobSqWm/GlscKGAMLB3yt39MU7E
USNkLKR3duA5jgoBE8VBjJagNcRGPnu86adMwD4os/7fSd3O4k7kwkyiVuGOrk27ipk7YPHEKQWz
+jtP1z7bGa7mMpwdnlawNV/Q3STpLXA+Hs1fXUR+hQQSLIJlKZQE9T8sX3GGbnkBT/x3bt9ad3tF
+M/oStuTIU2UybBinhU1eYEHIy+wpSxILLDLW9FwUUHP88fv0ZpnEEWi7WODmVVvX9WYoK0QFMPa
KjXviYAnIGLFfk7GNvp3pE/7VhfmqUs0Oi8H9c9w2UOLcSH1afOabvjCQF6x6KMx1q+bLj6YwJEJ
1AYfNx5vmvLatw604UecTFRqIOqqfc5NO/n0b7D3ENS1djg63To3hXFHD7sKhorI/dS/IWOOKXm0
sUSe9+OZKHP0jzTsgoJGZ/bnMIEIEFgAasXN8C9hlj/EZvCV9oKyXrsUhKsxR12ozzCtNGoitRly
Za8Hr4mABZOyau+hJpZcRSAqNn0nY6oRvAdifvreuxoGdQXigErAgTTyjlbaK40nLpRnugJRrgNl
X74v7oJrkreEsPJ7wCzHygS6kacQEmShx8565uz1uNVHnN1DXUoojjza1aDL2cQcGVb6yeSFvBv4
EQkMuHI9k9fboMYkegrqSxeTKTq3ssi97aB9Oal3BumW6KWYlDPphZNb6sUof5EDjqUk1w2G/5KK
ajkGUZwhCM2xQuxyKHefp1dqvRrBwJE/aZf1okdCPelxxyRqQtHou7EqSaOSwVW4uEqminZLUrtF
y/D3krIxA+td3qIBIzCre70DfIELcIgfGaq1sm7wO67WBsQpVgu14iaTtszYwv6f6XDiE1zBX27b
CkTZWzIqQQLpaWi8pza6Yuvw2Ydpem0NIQZTsKGhccVBAsmSKAbOjhAIEZf/96nY3jYgJQSBWCQd
2yE+2MlFDzktPm+BcF1t0FEtTkJMIqBdM1LYU6ZVTw2O5Wy2X6NFn2kAp32fsuCzqi2X5shGLnoX
wEnbiJvN71rVebT0tfdgQg2URsXPCa8oo/AAhxjo3k+P28/h94Vrf6pbBBpw+vP2orqUzDY5Wdpn
7LnZDgh6krKcnR/YcBPawNnOs7WnaE9Y2Z3GK3pOuQYI+0hxgtQsOgdHoHUP62Wg+gl7YxeEB5Zh
9ujBKeXONoj6zxkWDp2YDeLMhgZ9ZBEgPpb5V6IdpIzMlROKHXbqYv0bdWdSGRcF5x/sIeLDWZLL
k7GGyHL/nyHipkxFDJs+aXW6bhZPrd7ZzAQRPCJUNm0Y9KhxThT0uCQ4eDU0HGvdU1yZn/BcoPTt
NePOUstrhfGyga1snma77j+RFD8Hh2XKu0gT7EQLW4jNXYoloYrFJwsvaRxiYu4KQkOU6eMRtJKR
JAqifbq267TuICteE2GJmb59UcXQ0/uFhCJxa2WB4cxs6r/Fq3HkVuxY00WM83aiquyUvPdhRW8X
d8QuQFh60fcZL7deIlAZ8z3vDIu2J8mCmmkAuornEb+hsivhpCl5IoAJ0JpuqnvvBepPxmhU8NyS
AgIcf0veb7achgAsHYyWXwJrqlwDYK9JNLy94JhH0c6eDJgvtItZMd45+QAhMRCnoliKRhSfwvRM
NV1hB1MIf2w3sdzgp6eYgLMxaGNedyvNTBagBC7PStIbBKvdEsU5mYUPt86xKCrCMvStEMFtWw6k
tjIkhLe6baLvwjNTy6KShKBDfN7F7EXCrKcqz2ALVw9jTiMsFKkJJ0gcpnLxoMgCaMM0JGithK6G
U0JTtBjbQZWf7yWRKivStGcl3DtFahWYybK0AU+pXnbsM6n+e9M69+9OSJO+fOfubWLFMlxoseBn
2oP/Q7kZ/iVHpgIdW+xDp5r/xpZYgN0d7a/bMR+AnjCiic1Y6x083TumUeyeXZAPf8zk4MaRqu6K
4lIgeUlZvtqZmVqhEtmESsbfOALVnZ4V9K4WT6ZIPLSyDtouEiToiy2voK5XtB/x/4p537AIJQVb
65g3AQo2TflqEaK3Zr4EoRS5Hg5ux8LgZ+VUmm4OUlKcCGJWbWoQtbzMD89HPfgGNdXLTOLYJ299
zES1r8bfxgWdOi6CWy5YohH0mEhkBznxQb6xQPtimHJY5DY3Eq2S2hd+IuEQRtuCLCOvUmEiDOQM
ukAtSk+uWKDkWkyDWHHQHQUW83uAJE27k0N5ExyJY6uTIm6k1tDlydaZuxy07GomiLth0n8st2Yn
Y+wbh+9tt66eBEow6sepymdg91XjQP+hS6HhzUeofSgtg+ahW6E3mH+D1M6eVOW26AHMzMv78uEh
vu0UGekj7/tBDevr1G6w8Ps8apboyuD+MZByJx+fq0z40LhoO5Kdspl5TYmBIyc8nkVXmyl0gRVV
itxqld2FEy0+XNb7CAD0PPAb1fQFeZmHkpmMrm+noe6ZQ592pVVnxwmaHmDrAIDDRa+ITsS6XQBt
mjswigAmZWRk1wxXm93UzME15aXL8DKiJerLgM7BzViZmiBTMcDZnMLspnNvyX5NCesI3C46MnfB
uVpb9JT6lc14rb3JKrqk7RuePI++Q5uExhkTl8bv7FRcOyHtovs9g42uslhkXpF4+vrrUJyMvZ0M
8RWWD7K9yA1xpBcnM3czok21rG/sDVqx/LdiiM00KnWkI98Ih0wc1ouHPmhO0zrTNmfoIZ7iF7A0
ntLu+HK6t3dQ4a6Tqc74kxjJz7YZHwo4/Z9cxTnfAJsYL4SZZJeZH8ldoxUkvzKMgGu1TUvzCt0y
kYIYQ9Jyvc6v5/+/29ESqMBd/bFRG3WGLEGfNNvCgrd6Y6yotDDkilE3LJSJ4TWpaxxUyTQourpc
VyQvvPAuT+CclWPSZGW2fBcTK91qHJcTYzLvI5rhPnvWV9ZB1DgHQVxrkUof93KdqQcfqzjzlaW1
lHeqN06qu74VEYO4/3kCQcO1/YzM/s8ZzS95ulwBdGu8caURlZTZDN9m5XMB8iBAik04PpKtvcCI
q4l5noM4OOdta38BmrQuSj3bdAexEQF6EL3SjSbRTC1RSqP1jIiytVqUYEzJcLUAxz5BDFP8DJW8
PHivQvn10Wice9Ab+B6bj2h7buW6NsRt/RrUVmyzUoxb80gBneM9shpQG0fTFl0FL9vSfTEvH3au
gpcnvltfOfXbVa2FbvRRqTrrU4HZYJtKdTc8M/EBamo/nTsma0c7+6spvArnutdyhe00ES7CbbW/
oMuJdcvT8Qdt4d/+3TCPRL41CSsgUH+Jp3aIzu9ORG4wYSXTaZrmQS+LDAeVsgGIF9eR+Wx1fngP
ZZi+8xUYx166xOrSf8LYNp9Z9tev3UW2r85AVh9gqVEhJKTGn6XD1wMHr6QShAmRLoqbkUC4H98u
3rvEoSG0e/p+PDQj4veZE2KkKbfKv6T5MKT+svjBxJxGzh7t+Lf1eyt3Z0PkPT3kbv0pLzLr3345
8SB0inVoPH86Jz+sXyS9SWWRsBZJHooMNRrQ6rovFG9xn/JqtO255UU/RcQTlPOh7Kk3JZwIMNu7
V4LmIgkuRm/lrjYbDNPapGqeyd5qDojEvBTQmtqnMOhQuq7oxACb+Yyw5Xwf8Okz67YLzaSdY73L
5Xy7ylUdPVRgV50jyb4YJwSC9h0io3k+Ecfkv1CcBiyGcW2s1Ra9gtwbgUd4PPnzbQnz3UK4sadV
1yg2LLOCisHzVRc+JxhmhLqbyq7ofza2ceDhZxdDmwgUxh/e7r6NbDDTSH/LvAu0thAB5Qu2iwdi
9PBdpi8PCCeq//5URvhs1NTL9C+k4Oxz86oc3xO/k0iEE2QnwJqTlLDa+iqTfiHCT7yxSRxgzE1u
vLMCHaDb1okYnRCCspcVPkVVffZo3h5G+3Cc6qqLxw+/IJAviWEpHC2AFGF6ZkmkgpsLVQrwhMTC
2vkfNWGjzgZIsJHgIfrBpFMbSkCNe++wFJRhcYCbBjWfuDE9Av/tCPXSLgdPaXFs2N7/3HiGB1hI
vMZNbgi1Lf7V5n0qq/eYcKV/03tRDKzt2qegCKmInD/+1a9Q+XyypnQKlblgc0upbVSNrO2PzbUM
zxT2ue6TGKPTK8rmwnYRnLA0EslIKPpIhrKxcCcefDfBmOFNjV8D3p8Fsb6GkFtBwaFL3o7qwSP9
g0Tkvzpz0wgkPL2l5vkwDOZyFUImrzMjBAfdUXhf1pObEn7BX0A3YXlr6LWpYDm8A55Z91/HmMq8
+uHo8f+406+blxNneh44nQIqqISeqwC3zcClcJyTVQKpIzTS+OfaS9WtrrTK7dk7WgMkC5djAbkX
5ZSOD2tbZON/PmtmHnCoig+izZUoEceHpoCV9p9d1CvHDNdzAHM0q/BCOkNosv7i0dQeTD4yUmze
ou5orqOmB61y0G4KjnnzHCr4cxJOwkH5WF+TUOxRLkYkVi8PWWdyfSGvIdTRtRE3zhTi3OCmjWrY
fXwpb/aId9litautnI0BPx3WlECRVDrlB3knvdLnPVTTPMVMr6AHrVAcfML2gbbr941eUhiSkWmL
hjd2OD4Mf0kLPmwdoPMtBx4af/EXskVI6NFUvvtsJEB4S3QL4BvX8KZM2/RY8gBjLOGKyPjx24dA
HaAMZOb20yu1lndZ+W71FRDMjuRBVNtNWes7O3klHKkDymbyc2jRTJAD7Ipr20kWW9mc8OwbiLu2
9OkP48Prfdsz9PRUkcSB0wKnRwsiP3VvKyfaGBfVuCWM/idULbly3f5pkwnIhmrhjWOenMPve27H
nx5UkJWtCdj08lqzYGxBP5XCxiHko+hkejapGVxdxF9Y6D4rFUEQoyLDSE/gODqkIFzk7FySOc02
q7nN1m2iHtnxnc/S8yl9rPpoqgrL6tRVUWZASUyVTlbeEkTa0q2k7PJJr2qm2SjFOWcN44U+IZB4
Q11nxnOFnld98H5tDWmz0ldgcveHTvb6D0VyG549qs+qHv4bS2NP+DCQKINGnOzAzVs/jD4E+WkW
8FAhjGlfsF0/E6xc/G5lpRKhq8M8m+Yptz7z39A4NYm6NV81P/xk/nPwg8UOarggacBw7zeLYXP6
E6NS5yFrD9jrUrQam6PE3DsIl7/V2T+ugglfOHyc/v4uhZw1HqzFIlpockJVv/Fi44dzyeW/I8im
aPkSENDDCmWbT9L7JuYdAK7sbJWMLgOgCu7Hftz65FR6X4oEm6e/Fecnae8pFF3vE3zR7P1EVQIa
GeTj+uszj3KhWRTRVjZgyDMPYX+s0Si8b3CyJSxw6waHI/TxfQW0EjMfhvdNwrAleWKy1RM1iasX
xebKQiJG06lzThGBZZ+YPBseZOu1pxQj+HMyPphtg5ygalxiPx4hxq5kQT4Wc0QQOwBZBCLQpA/i
ytccByYC8mSyXDDKt/nnCCdXrkUi6pbg4RfOWMz9bNDHBfSwevMUvn92WTEQSGl3ABc7caS3Bu1u
FFeAf7nUt+/KmxnPU1UDoV6RXtN5ACKur4/IEG7g+ZtZs18l1SMv5CDHEjp8wz3UkTXT9Ht2e0v0
j0Avk4S8hF6hgGO3SBdztQ7F3fmgFeKMKTEkHZdYhdYlIBsyB9PgC5OhHU5CvUg/EcrDbLGmQTcf
KD8Ed3mcvD7/R3IdTT0BanlBAQWSN6ZwaxC6IxzSYf38eFzDEC3QR6x5AVG0UMssuOfQXAsVM96o
Kt/lrgs1VMUln0wendDK8rfHRNmhlW48Wz8KFOs1wLaI2UV1uOWg7RYNYK2fG7LiTyMqozD1K96+
xZaijYRdGleH/mHP/uIVvekeloWGwRU9BBN6zOWapYvI94IfYq4aGkq8JsYDCSVhmv40qHAH/i4P
cf/Z0iiQ6dXbMY5ktB5jDpxreVRAxH/I1Tu1XhIBf5FgN5tUIMuqzubDXbHkp4rg6h0OJGNi8u/3
4WBgy4jVTFfvvyyAsxktIGP4bg1CHAEAotxKzA3rvxnmR63zesWewUuix40sa5/K/mbEquMX3bGy
47Uk+8jd1DgpnnpmoQDMZodTQbDd+Pgf22qn0sjdBFsl0/O00ibJddox+abwvnSrgazggNYCa1NE
1YdKEldLipg/LV0nCP8OKnnCNDamJH3681UfSqnjSfkBGmzWxUU83F+nfGYIQFslJJBuh/RGygLh
LY7Uw3IqF1ZqCltJcayhO/rxw1vNYOY1zMRrYf+ZIxh7iB/9DsuDS4Rzj0d6DGOKbCKqVy/qI/eX
hAoKxrc0FbBcE41b7Wrl1FSM1VKdyMdtoJUWUrfdP6xY7D38Al32i0ns+IAi7b22vX8R5oH270pa
bzfU//1EqKwL1Lf3cQ1M7gKmNbjvf95ebTB+OwhVRg3KeGDx/EajHmVGL69m871skSfQzI2Vb5ez
2DP54W4nd8dwMzwQ+hZ94nAezkWcsoy8n60S5wQrjao4tkQuEuS+4W9SpPwSSKzXXCRY2hcVNOKm
ZWLYm52srNOKt48gnLsk6+plZ0k3KawDIlxS7d5AOR+uwFUoXNEbKnh3trnZ0H6vgdJkM/wxErDU
/OhNo4pj9iQqWy31DlbPkAJXnJDAbPIzmj8padJPXZRmEQXguVjuUXRwJVVaPQGR+HwEpNICoCcz
LPxK4A6Y0yOavS4gfUCjx2UqM8wVvMAH9QOm9+bWRYeUQ4cu/KcQvSjiA2hIQN0AHwlYVk9cuFJG
k56dVeHJWLGQHyZsSyEhkCiEH4sTUxy5Z66sboNpowzlqJZzohKeQvJz8FUd6q2S9g4zFLzyaKJl
p7nJw53ZAmf3wBi8cyRQMLQOoxRqNGZjmqChK2TRDd8UL+aL/PDHRYWO/lcYzQOslInh+5B/Or38
Xyb32Lo98Oowy1eFVqr/Gf6HoShny1k2oZH4Rhoh0PYvY85A5RXCIRdmEDP8RVUA36J/ZJLZxSKB
f28m2gn0RSHndvAakxhzgtrHXFqpfQnH/yB2OoUo5Fv5MkM65bv0C0H1ljvt+tTKN3i8ZU9T9yLl
vkh8YL+6A8cAc/ira90SfDmyXQduTJBs1OOwyzTAKq3drRbC4jeBJ/qrVFPIZODZVhwO1L6gKm9H
iJDAB75fbT7Or2tE3Eoh5mnFBy1V8NygnvohESu2v39X3nWxvcXRBqMTgt1j3UeQ7Xm+BHpH3XXt
kFpaxawZJVRepiK9CZew/5FsaS+lnPcz6NrjkBvCAD176yB2B81WIEpwDJuZQsdW5MCUxeK2D1vp
anvOhT0dtLtpheO3yj7+3RgPXzKae+EZsKzhvgOeJFelR5xfuzlLvcwhjr8CKphL0fbxO0KTApnw
DuRbi5z2/nZQ3xCXAqxYuH8iVikrQJYTXjTpPDz3BxWG4PUrYLol5vIXIYW/tIEn7hZxE/mHpY5d
D8/1tan4rX3arQOZVdDAXMgd9p/vD++G1QzayocwcoNpCDGRNEOJytmQg8IhXC0tK3oJ0MT3fY4g
dgIByAEaeUkO0bZzifyUiO9G2UNLTxpOBXYhr5zvN2MdYxFxqAiJnvC4KL7efyl1ih816rKu1Ahz
qeeCFeVH8MaWDdjfdiQgdzwOanuhmy4ee7XAm4jcof3VUVc3SYWKV/KaHFqOhYnz3/JQFc/voSm/
xONB26UaE1YVXwDpcyIKqraIzh7tvHGtZd9NDEucVyG/ObTLWiesfLxYdK9MRa0aMRVTvw7NqaWE
Ci57mtnvGfY3MQLGDjWZqtOSLm1a0Rym31UHz/CcpPGXsSwfVe4uK1F6NS7ijY+Y/Vz/2oTBva9A
I5tExnRu6M4tvJTloHuG5QMKozE+md1eOXnqKUS/YsdMcK8GtmyLqnW0G+QcRhHuBIpi7rE3759s
aHLA0MpIzEdeHdWWFl9OQJX57KSCR1HCmeHv9kgEmYeFKC5wolnmxewQIz6lskygIryNjY/sCFV8
CZeAkgQjSyF3wSOoK6eqKBD6b0wyKJJkSMCv7WYi0GVrhWyndyAQflSJYMyQEXCZDT5TEpyJaX7V
v+deBB0Qh9TqaNI3J4VEJyG3yZy4Wa5dtd8u0E8MfMpWWU4olmc75Edxf+hbxoI8VVNXl71Dyv+M
zCkOd/pEYmOO1v6oTVM6hic1KfJ3LWgpub3DABL1lnaUxf3XZJ2Kf+z//alT45Ii5kTMFJtgim8p
Y3oR85NMVjjlVk7ML9SV9njcqEcTanH7utoIyVElBcoSUTw3WGXJ38ZdTIihjWl+ZispgnQqDbY5
cmy8qVL/PnXlmhJt1EcsS7bcO/a8D6eqS5fgB5MR44Atir1SdaVXAQZX2Lp4ITUZe9P1TIApZe82
FE5QFEjb3S9pSUqjYjvox7obeas0U1l4LB+ef/ZazXVBn77n2cXzDNyjVhF2HCPF72JjsyB45AKC
h7nreG+Juq0P2t4ortjB1SIjsBmQTsJW0n8iBOEiTgq7oe067z/KAekENXh4+iWeCi30OzVimOH4
DiPgDSs53wsKAl75P43VNnE4o4ffPOkA3MNv/qY4jmtz5w99eKkygUBuz+G6euEmYsr6qC/wi9T3
rjjxAkWAa/WMyp4pvkoBSmZhasC+pX8xkXhOlL9TIOOpJkOJIvw72DG5bmPZaDyJ45dE+w4Z7mju
afbdPwnvubVT963o1WtOtsxgNHYG2pm0BFEDurQHugI8gUnxlSRdPoq4c8su/2964qNmhFBHVtZ1
qEnzIGXmfWss4RDVvNPDtbu06vHq36wTvf4PyVhpB+BHyU7R6hARjimcN1vB3B9ZbpYR2v+JRGxP
5Zih7KNtgtf1m+mVS4gzzCGO1UbHuVZa9CKCF64q1W4EyjiwVbKnT4TNhqroqjO6wJFUAsKDTpi3
6QRRtQ2jIFDl4xuvpXhdXiRiPIvhEEWuKzOwB9NuhNNleCFOTVkpcCRms78SFUnIy5uUMTVNCkI2
l7ZZdOOvITwaSOaMKl5VgwS2O3ZXc9bYOoh1xWn3dU0qBvOSdei1IMhZT6XRZVqkItFCVuJdDKcm
KUT4vhiOG6fgfe1ZYGfx7z5yit/MtxlLxBOla8jK77nel9pK+1wO4T/Wx/WdAi9BDHpjdZMi3XgE
/YCCszVsTDY/K7ImibWgOhn+KR3rPAtPDAlTKmcByKGDLEJrkqI0LlTgPY1vZX6zZyvrWixloSfs
65LXVBYFsy9cv6suVfld2nsW5GocN1fSWybmUqJZO8qOGfkq5S8yvfMLi5liTRPxsWHB8N6aT846
PxdTJPRr3dnc8kCm9mB+EJB9CQze7wuJqJOGnTgEVrUhbLTQUPF1UChm+pUjl76+xNQOYCfphfqU
JIeeHjylJmSNNErqNxD1aaoja5YkWO4a9o7mTcoVHy+/P80qscy0ZBLpA9i6gY2ltKGla/x6pR4C
uMsIWtdMuR8bzCNbg3D3IspFuIf6CD+J4f0+oJo3DMpE1meEplkqQr7s+tB0ioh6A3JJr4ZmKsVf
3FgwMcgHBPk8eYxacndpmBQPswGTE72wu0zU2gPxKtrXN/8TQHusE5wNZMwXTXAMmv6Il66Ulqc5
vM32z36rhNva++Ge6BkCuU4qXmqYzbV0mfOVlaQzgC5EX20NYsSCz6RVykmMaWFoTQyGOB+wyxkA
Pnzy5S5UbisCa2l158d1VqvfLUi1Myap+p4GBbHpemXmIn3uaJscPDd07nB+CknxCox7OOvZjAjo
xqt/ErRPQ0/MKfnzjB9mnp86kToGPn58cayUZoIx5ExTPzZ5G3BEQ1WJpOp7w1Zva+of+1/v473S
HjWpxGBI7zhLt7y3lw2DIhn7vB3BtCr6REVrxY2YDqMw0b5njObf8CfgOdFYKg1Cq4TBNKNexm4G
3vJ+pJOOJvRFugSSJBZaCHTvDrMVyqquIYJcndQCfwHRXOPxxsze2x4uI2Yt3Oglh/pRQQoLEbX6
xXYokOiTsSCPF1+hV0qWb8IM/byUyrAI5bZhjx+6qb/PsuMAiSLUazhW/3EzYFCrx+CI4Q2trOc3
++YE22pQg0nPBlQzC/DBX2MLzBefu9x32ahccZ9/yb52ug7gWtCGhM0R3iHt/o2jK2oIpAPKPQHD
b9HfYYh8MuE+XfqFyEnToktt9lp2IlEXKZH0sF254f+k+qVvi/J1q5nUITK7/9Axbz5X/ZyeqCvx
VvNFEcT92aMYpXJ32IMOz8tVo5Wq1ZVVsJhdyAwORFTAkWpFIwLmuH088NV2kCgerEf4z3BHX+xb
pYsY7c7kckPa3wAsMiNrkvCCXnPKaWPsC1plEJdd4qN9dcD8QFhvAlnvxby3jPgQ+eGMznwGEaMv
UHjS/Ni9cAl8xaqz1GSB9O5CCKSOaCVVeOO+XmI5o7OKy8pbT36atnz0Wz5tIEH4WR2RYAq0iV0+
480zaWQG+si8A/VALYA/PhVqTMPMjcwk744U+eXAq96Fq2MKIcO/59d7h4OWmarVrz9gn3fMyMVh
Ya2p+j1El4hyRIF9x1EO9ZRMeoycpInFgk3CAqBOU/2BtETfIenl49vFbRG/Og/OVwLaMXYO20hZ
YywuhlZtmSi1WAxUT9syDdDebN8hiphkYiZ+LrwP2TjWy0SaOqCuY0biP4yUqq5VimKDyI0yUcdf
xPm8qtI0JAF7oJuVyAQlV3l+Z5d1c5G+ep9hITXdAApX0S9xkssSxc8el17QSLkPXBWqyW1IRsfy
Yc7TeYEh5DjWPeIryq5zR+eyEVVUKlpgrnpggkgBhpGPwFl6Xj2Y8jhaYFKCxG5dYOu3D3TGfT4r
UV9uxS4cFVr75pqxbdgDnUKc36JSjGGW++sXEZjHXXlWcCcSKkIBPVzdCwgX+hDrJagzkk2cW7Gx
zKj8PwCaLZH16Eo9S1EQwwjVmMXkpyZDbKYJwspnRpLnAma5wZ5HtcX0W8CikXlivzKPjClTYfoU
FQ20rnrDfhaa1BeI2zdOeK719VJoe7SmYOvB13CQY+SZMT6ynOE6MKkZ5oI4RLGcmfHcrhKEil1f
PPh4h79sDNXI2TmvJeE3inp3rzM/brz34eoy2DO1D2eKAMA4w1rbVu2Lk+ouvpvQO3JBU3C9HE8H
ZDTP0y5qAUaePL8zHxfZR09AZ0qHfnKgWdIBLnJaKjTlnmnhs3DWcJ3tGrRxJOBUCpKtPCk6ixE2
lZIDud+SM89NgjZhFZdSm7Dm1w6Tdzquf6MYk9W0np5AQk1BOOPxMnbyzjf/9Rj3qDsWGKEU+7sx
sHVSf/WU8XG8yKN1CEAXp6z8SN0Xlc1oX0ri9tJQl9zW3TPFyfuvU3++xQ6mSEPnUpMjpHSxieRl
m/6Rapm0RfLw3RRqd5V7uRXIXA2sDbuveW7pkFkgZg2ClOEaFJnbrzjR/CQQnB8fg5iJtJ2CZgCV
FgmR6KFzuUXUvtWA7+Ta/1dE4CMaSbkM1F7nsSFukw8QHZ9hqMTJivmUO5/YUBQ4hVmrCILF0U35
l5eQGRKhvsa3EXH6xuSQuhkfd6eJPzK7NHoOdxTFzyqHNWzNF6V6c0iCW07dyRRTAM8xkXgPWdLq
WNTqZa/6D76UYr25SXWEA1oJpfvRddZBXlIj0KqqYKchjl09SQ4oiOWRRAmg0u5+vrdYnIYFbjNA
HvtCrHgvjSWfFO3aMJaRYgxtsTP0cbX0kXgIqg/iRM18cEoTOUnmloAGrfPKxBBZ8Tp9B1RV6rj1
5trSwyrPeWcZMi4Z7I79rk5YcCX7VFM2EMvci9dMjmCq0+j0Erox2otLwTNzrivHAyAeJSB08th+
XLLn1YCXtIam5ijkV1y/Z8S9bRtJ32+R0Ny3Kh4e+MkSVif1Qq3H6l5YYU7E5j4MTbBG4/zV3MJy
Dfukm9yEPM/XfBzQUYjvifWQ8FcwJk6O7W8CzH8kkxBJRZ5vS771R/kfksabGgtkjCi06p7sll8s
XHEl2l90qYXhcwJZTNK4DtIzz2n+9ffMNG4LVTjaT9WlaFhSZtQhf5odeh7Wg6xcKFX6jxTBLQuy
Ka3Io/PdOcwFYjl+TNt8vHqBerCzolG/QAtfPIxGUXEM/PnPAkHEGdDBkQ6C85QGKV7lX5ZWId8g
tnc7BLP8gXUDpI5F77EYCh0wr846sSQWHD9eQrdxM1kScgiPFk0LacpHMydu7J03I5hBWTvIGlyS
jv/VPpEMX2QifGEtqpIo951rDOztrmmr1OTvskOhQwJNFJT2JpCUc9dDAZlhr2yqRVqdtFqkn+/K
ONVueUIdGbqBgyLmKbkMiCB5qlwKPzRJWBOxXDHYmzbnCYbgNukNHJD4R6my7hLn+uCV2aMbhMqs
Uy7RTbEH1kkF/sDDYRjBBbR22L/+RryZmahFoG+VdOa/YR7xsRApOw9LOuUC0lzkovTyDYnjcSI/
h1XwdVxcRpw+GxLWj32bdR0PhqdoNVV+ZSrp5UuaLMP5sY6I8Nl+6iMiULNkeZgeYz7LAuBbWdTJ
OtEDmBIB8srQawoa+GkRwSw1txZUD2SlfcizNILjKFKjWZLyZBIdQ1TghtuWDlHoporB9Q07/cVg
cWeOz3H1KpS2F6mHeE0nmBMvSUvocjkvkq1hwuuVst7e5ZBpwQ2p01bi2ZW1tMNils8N1RIh7hVh
vUNYGqqcyxW27+5mPkofNRBpac5wJeNXE8jAOla3Xahg/CZTxIHjgM1RzK+ZVQHIbKfrj7DVVGf6
q1bJyq4w19tDyy7t5ozOEtPDUypZsdt/6pQz7EgS/3eF35XYNSb2d1WkOgmlyXHXDGM0mATCtlwU
++hY04PGO85rlFECZfCuBN6Zbk4qhhOsdfpJl1BVlwJuPuJcYGAP7qV6gFEDrV1/IPn5wrZ32mIQ
dPWh5XQdILpJgF8yYuB3Kd/qj833npfgFAtIBxBqatZFFN2WNvO2tHw2CL6rXXjxj581p/Jo3ydM
PjDc3EN+HyPHghf9E9azlSTi8GLhdvVSRJJj0lT00rgp/3gm0Hr4qL8UFBrNpTHV34JUn6e4jjuX
l4lt+aBU6/fJDNQrMA/F8QNMV2ddfn34b/fzH/n+amHPte81zIZA4DHv7V6f19wCE2cI1D4JLVlm
SGCAPAz2D7TS6Si+eS5aotczr7h68peKsf1yRiCWshbemZHNyI4qTIxESM9Z/IYBbOVZbI49ih1f
UBGuj2Qby3J9iisz6lpEmptY8VZEr2cUWJTgZxgOV0LdgpR3YUHfqAHgW5MrUmSYobCQfiNdSKiQ
kSAfxPs0kX6ZF5gPGudNOakVBTUoxgLavfE7mlL1FMdMlHRU5oI5iRUQ5X8LUzT+H8GINx7OwWhP
c4KsmqJccC7E4yjkojcu4Mg5sBE6Scnz4lnwMDIIqtcfGEn/tCFG1k4fhL73Fwhtdn+AR/B5xR66
MCe1wdA+Fv4JqG5cU7YrLjnfRJYZmF3xSj/1arzePopSKL3XWs8n8BrR4zY0/lYKRXtt301v6Z2P
MPTFueNXRZBGyllkVL89q/GEKbTLRrvp049/p7+CQhW4lnyWi2pN88l3lu/t49NG1wQOOeCzO+Zv
JuqXpGURf9FwRB5/796kkymkQK1TPzwelB4IevulRwJYlX1zND2ggrhaABjgu2YF6VAy+lSlnd6V
jbTBbUk0XMrYpypYqm1zBmRbUuK3sKUP1nqpdTbn+ndhkhNHaMfjlBLmOt2rdpRdV2VvRHlv83Mo
v4gpFF5bCnEeqio7c20conGjsjrqyYyjDV/klPCDZ2peVp0kHet1kak874e6FnB0gK1JHqQ7UKlc
92QKGJMs8SvUNj/Dp4tCh19jnwjp4iYj9dZeHitWjN6inDCH8tE9OLfZlUbnUFZbr2sy2oSja6ea
NjN9f8UtTyQHoiUZX/VXAlKaWKLeHko6kd7V6ccMHBgLtl0CiC0XMSd7/m9rckUY1DBSV0uzsMN7
Y6bjNYlIfsHXEnQFL/Z7sX6dcUWet8JBzQlOOibrm1p9PNn5+0B/3SVZ8m5yW+jSHnr8N7WrGnK8
vyj0QvdfV0HSSV9ZjqBn8O6l1GHHNg1dMy4b3Vk9VtNwxmN64qEpdKGDv5d8noUiXDSU+S+q83IF
ZN6e4B8I5BHDbLMRpMqp8Fq4aGIXkilPUjTX6kZN75XorrvcSo+8n+xrZzjX471zbHPk5pZ/Au/P
Ek1HuSZkvI+McTgjOZGotcLVysYHhT8XxwUwdZLUYlXxNLT6ytQXHyNFkLaUK/QJGc0uyHgJWjsm
qGcVDjgPUUgUSiyCsBdlEHWLd0dFWveaqMt47wZRDSXShv9TmcaF2yDZXcQ1RlqF2RUBbai2t8Kc
fTjtRv1rMCb2scA06e417Y+rFVBWZgUeWsPX0bXvNSOtjkC8HxBiVFTOsvb1XcC7Rb7SURWrKf1i
DlLSxjO3gZZdw58N2RoHzG/ZwlKRqnLR345umw0J2gBTPzLzw0Uhg5IWAGCQ0I60hHOzfNzVOl6Q
7Z3YClXgw/OGw62JaBzX0+SWeX3k4N/82jzc7uyoheGpUscOHnLk2werBuzOfsjXNNIt7BmwOelb
uA/+ndBinPN6n0Fw7kGJSyhN83SxcWz7nJgQYJEoAS89tqf7bgo2FvGlZvMLDiR7hiDb/4xSWXim
uecuTEZUt2aJp1iJJbHm4NjvcPSvcJaM/Xr4dui8kCQRNRYykH1gE+MRVySByQQkQQ1uoDhuPLRk
eLP9/DPeXGOtjD58IBXdv8t4DJvMZpAR4d2SU1mfhfrgQr7B0YYpvVG3OQU3kMC9UQVRTIM7x7ta
/Nk++qX/X0K5jRigrkXc63TLiGAdt/iEPJfm5BuENlZ1QAFskgVJfZD96tKw78zGqIBe/J36q5n/
OSZbnbf/1DZ3X2U+E/50H+mqvXHbjku1G2U7ORvpWRpaAq2kygn4N2a/Jxfzx9uY3U+neofpzmuL
dZitpJUzdsUUFjJjhCLTITlanOv4lS+sMHxAH6mhADrNDTTNGwMKLcrwBWPOj01LT62krHU5+ZlU
cWhVXe11/iDg7uOM2xHr/TWLokuCAtYhY9aRBOUWp0NqAzOXAWkgcsGW0UEDGKH7duFvF6adR5eW
SMyjFrjPiptRZomah4P2XOAuGRyIFoOdgzrjBBm0qdukje4oO/4xA9uL/pVyoHQUvDDXVwdkTmK8
eJRYX+MIATFOND4u6pRbEAtYYRb1b7myfbSSLXE8mr+rY7FLHAAhS1NFF5ayBmi1mVQsr1lJNxF0
CKvUi+b4E4SWdDeZgVQFJAQ1tH+CbiR46TaCDztDdFNZGzO05xEmxhWofdxxK4cEC2FxH8/DbEB4
ztnCr6u3CdYGT/yWor0PeSq8PRYtOkN5LNxsstVMsN/ooYwYbuaaZ6RyrGJlU2fazZiwzZ5SI+0s
f+8sftJdzqE9Joaiw8od1o9yvnHr0vUl3roBg+yVrPnxc2ieGBTfzISnM2UwUuZt2TsbFgrfrXXi
h4K7cBXeGkL+4AsSMTBmbP1YvgliD+mCRm2YKJkmMtFCW9DpEhWsrjgqoKisRb24ijRoZD8Hce9O
9X/27E4Xb4GKcoTBjmHCii7COrGHSOxQ3Q6/1rRvqQkIb7gQP/XkNDB98x+MI8rjz/ucJjGLhtdb
6t6vMQz/p6SXMm0umJ+cX1k6jqJj1ToTi8zclThMsh2EqCTHDX6txeChb/6QiIbuzBS1zr7xM4zB
Fyx2XdRZCvj7C3V1HBd5Safzgk4dHLHpzfwaTxTquE9C8ekW5MZ0BzLvEozpgbFgz1bh414rNBGC
Diz/6IAloHLhT3RPKYueL/3t+eU7u88AqtYhf9VyFwi22BjuFY1TC5SRJtXshbZs0x5T+im43aBs
daCYgynRC4MIA8QWylPb51F4WiWU2xjQhGZ+U+wUUHaYG7wLUDBALqlWe8WLReQZLIiCAc58h82i
XPZgfLrxSZZDBWFDuS/aFRkYR82dNOS0Nhi8go7tML328B/59d8rOje5syvZhjmzrudSdFYVL/+T
Y+f1h27q59zR66nbu8VW8lyFdOIzPciHY6/eedOb3vqWpqWi/wwNPFFkeAY07ej5CiR1h3qdmUAf
fAscV96iOqswTP6TSBZ1H6PP9VQ+wDWW0WfUT6HLYgyU1/PzpdBoWBRLi3ShIZMz5jh1bVObHZ54
uiqivs1SzBhO+O5qzDrY+CnK1cxevr/0nz2X28X8HZwVXcrV9714JNppQqrAZ13yoS7P/XWLJ0hr
hPUK+pQbR+iiGMQ0KBqJcRn6CgZRNDzN1tsoTTjgA2b/KC+RO5KwIi5FWOETC0TJgCCBDSl2jcpt
lpofG1HMp2MX3FNVllc/smP1a2zZdF4hcUR2ixW+WFAvRwiK2Ehh+Dybz0btCktMhtoQfxMYd0/G
/h2KD+owZTpnU4R1xiQIRnb5xQuqq8j6FYQ2iv05Mfq6+PeCufIUbPrQoHCX2GxeWewbVGQLjnfn
nFxmOLnWUDkuq19NTfWLxVkgQcy4ZeHSif7x/T9Ync22u+JoMEGN1GnYAQxb1WD9rvR3e/d9VYYW
bEZupCvo5dYR1UYcZjkbnlcD233plUj/tOR36bYvdB7x1x6zN46C0dW2P1Lvbj+jvwADo4W/kcIE
e7my7A0p4GVhLwJurkfphFJm40ygPAftx0mCVXYT6uA46ZLHs890xja6cRSrHbONaxMNIm1Ald++
E8YFCV+0uo+vBr5BrlblwxQ9FVAKnycEQSHOha7/djfcP9cA/NszRlXEQ1QzewNudBw9eYaFxRDV
1NMgWhj9mmYq/ZZiJuZ6SpkaGh/W1X6d3pVnRfqMau0IiOrJcViuQuKXoKBv/igkXwupkTSZbdNM
XI1iWXORJUM89NlkP2BWnMEqh6Pg/D1KaSvT+wxhAY9WpXEOZ3Ew3E1SRhhjOj1ENGn8+Vm66ZcY
uP/VI8mA5zQW1WuEniaJkDmMiWZdh/HstD9dOUXliDTcWQqZQUD2OSj4DAUjBz0tXofpx1aXTB0P
dRdJdyB1OCU9JLrSZeunvv3IsZEJgZBDzwkp6nzk6vaxAJ3A5iDyDtWsKsou9QYfWqWxUkY4GcCc
mJHfvvRzoCAow3K7aRCfldaUq7Nccz8G4BrBSvM4ik5+Zt1MwdxMVMTat0D5iMBw2TIvDiZUx+8o
4CTWw4EYUX41kJu+1eg3DXfwPTn04FJmZQxPw6ao76Rymm8u36D2OdBvwTXubboKDzCZ88llnEVS
FqnSMQOJjjZRUYnv54aLyR2eNWfLUWi2KhbCgPpGy3FjGgEnTnqJ8vVnxu71NvsujlREcROXdmLE
zQu3N70hB5+5ldkcCXUUwfxoLsLunKgO4Pz85zUnpwVK100k1F/Bz6H9sAkFOiZFf7xOwUblNg8v
CsLKqz9ElOXxiTUWR5r9j7zV4ajKKystKx8twjtQdacpHZUgcPB5NieH8Uw76IXwrsk/Oh2ItF7b
F/f7Hw6Zfq66APWhJ0riZXBPUR5nSlzppUHF/BrlLKh+LKEjRzquOOlkHzttj5RqqoKwx470l1ro
pli+Bvv3kfwGQvv2uVJfy2G2K0Nj8JelB8K1JIDLbl6v3mSiEhEBjMTHOD2K9kmoabjnW9wMA6J+
vIAYujqITzBZ3z3+UnBZJXtWNAx/7teQpBY8G93sp4DEO5K8Zl6dnRFad4cMDAK/RiuDqlRN1YxI
YCnBYxQmIwNzhBMA2AXy7TFrlkFJo4aIIR+oCAOt4M+r3A5pa/aAzLIBk0ZwxDFQAcYEgOdJc1EL
HS7y1PZ8ben35ymb3SjqXzcbl56qH/NM2VzXKIr61g6RREbjgvSr7cCmdj4OGcMUWxCSjg5nu2Q0
9eJ4riALwJ16/mTRs/0fBOD4Jmi3ys67eKxerPhhgrzGKPqI3zqrXRn6g8RkfATbQcc7rI5jL1w5
AOUa4Q06KeTZuJmDbGWgfOcAoN1g764bmKyJFBh3Vv9sI/4TUINABIHbWudUzKEsvGhyBrpDCrBW
3SqprBi/5qmd58Os3IofIdl4RcZuY7ewuP4hHXZctTsqOeTfnftnJfJ81uuJeY8jPC4w3kMeFgr3
JilYtFuLhObMYJeXvzfEy6I3Kp81CNhw6dPJlqOFeB0GwmEhrKqMiwlU8hAxo1PRuTdQ+aTvwHYL
iAB1IgQ7rPJNkXR1wD7H5/od6h63+FXeByDCTkM7Je+EvBI2WtXc9oZQCQ3xpw3kMHDVnyC0uzRq
oS8JcZnsdImP3rwWJWnez7WwgdLjFKjXIF6cJVAjdnWceKcvxPb58MyFd6+Yv+daviEO/JWeigCT
fBCY2p8Dy7VlEpReA8BUS6WiVDdrsooC/NxzQtIY8iTVQtjH0mXGOlsNlFNDXgUB7EuIst4C5phN
e7lr5KP4aZRXekbF9SGpk29NH0B4ngh5N12anQf8lJwDnRXK0qbcdCFcVX2N4HxASRqWtbHdAGU+
Smcg/j2cWNAm7Y0/8qveoKYro9H0A7jyzoKX/wXVf80qQdwjreKOKdKeIYM1Mn/OnE8a3x2ToWdH
gRL3cNbdY4M7tDbn5y59x59OvWTswOb4fEyZMBVaistqsEgrIc0YmQ1w03BbSWqZBYFQDOqxHHZ1
7F+82/FlgZxrJ3VvyPHqQRuMjVNRQdIb5wZCIsS30/9yKo2K6VjApDEsbNW6SE2F011UoUa4I1sh
/EyO3ojL4DDjP+9Q3GqByqrf8eYWAj/7CQkI4uSmpdjWHca4ajzaxcyKFCiXCcuXDBy2Y7YHNtAT
TIEI74sq3pacf1MKD1Gzl5btt0hGzE5vDzXeXPZWejdmCyG/vfNLj3DrMq6bVbryuzoQQIlnFM71
2iTSLPSP6+2MMUy2/7A0gMwVegAqXxG/gHkMkv1Uf75z+ii0iUHZua8Sd4N4aJp7eMwZUx1hdSi4
QBL6F0dfzskjCeVhxwNpBXanFMlP248l/Ug9UYzoQJQCOcnUGHvXHZOYoR9uhNHBCI23Hmsj+VcK
1TwYdAdqE9inSEln/9PIVrvvCXvybRSBoJw8OdilYkd9i0y9whEXmfHAMai9bJ4WpUA95qsZZ3uP
ZO+TFDkXWjTyLnx7Bz7tUCBZXSGO+fkoFltr8N5Dsp5bFDbhs2MTqn/QDThiVj6c6+7NwpmrAToh
+IcjRWqrwLT5Nguvbh+kYr52Auzz4jxRdz2PBiUPhY++j90omK5J+mICmzBNKiWtAk5MRBYwnv5R
lE9hF/A1VM/TGrthdq36GfNKcRDjTs/NvCz0DM683fAwk/Rr5kjQNzhScvkBBpmrIHUq7+mXrIOY
8aMhkVkl2z7Wx41aw+UMjTUZmQyEmC18o0Q7zCJ45TLtzxQVmJYdbfz2G94Vgi6Odl5DAcwcD0ci
XXL/5SvXPN7duKCTV6T8/22cfXcKd0h8xBP7cMn03xND+9VczlcmCThF8gNcVl8TYXij6i7SHOOC
uqpNqK5sjNQaSJ5z6O8r1y0Gd4bsEGJ0YHMQzFy0VAqwNeiCcxUlVjxUVtX/oLrLrkDEguXOHQmz
XharEnGSDbzg/LKJa8s/idyHqFaTKjWQysJ6AbzyERjWun7tY/NdKlJY1jvflclMw+v8kK4MIAfU
bEUIyDrI0YoigKVfPs3xCsx1fka3u/0AMRTCjkhi4fQnW+gd+YCyIVYVjnSbTxpLR/Ekyc5de4am
0Vd28GJMLWW9dOs1/qEOYOyKJLRNkyZbCPkp2cW5lKxSkJcySYB9ZQfgBoC4//izarFmU7DKi/+v
H4/A+XqUPSsPLuzkRFf7DrFBssXPySexpU5UwjdLyXFkIgIZgHuvhg6iLf3iZKcZKYroKlpeOEcH
EC1wLFb4SLQ0BZcx7MWrS+ZGmqJXBXl3UVlPUA96PBszlUJa2kqttbInqtfniq9+rIZ8pithEqbw
Hn74f+xmu7oHmHOjFznnojuJkXWRqJS15hbvouysS+7pb656+qTttI0JUQrKo1Qt7lqCXPuIN9yy
gduIITvOz2WmucLUD2PEOYcyZ8VohtfDkns+oX71FN7bZbwzMcXgkRFh9H3Wjmw5Yq70fbrAgjPG
g6WDzQ+PAoIsKtqijIIHhQgFEXxysqNIS86tqKnloUAzMdhVw4tdLLSdueahYb+hbNdu2Z9FJAQs
ZjWBmjmUmRSAFlhKIFJcaDTKDjvCu8UYOiep4LLyn8+QMlt2AaM4wQ7Kx5A/x0XzM1A6/54Xubk3
0TZ8kW5FiccN7YLlNtNo61Ld+Ig79+y7KR5yhT0Z4jjd3IBLgdTzLG/JZaKkk4qMy9qS+LqYMZ4+
2O0xRFzbrjD8YqTs84bw105+FnOYe2VcsaKEvyJi25ZPQJ8G2ekx4LN7jb9IbFjSOJg9sqLrVnSo
pWa4+1tsZbyrf9Gs0aNloU/MjnMT5aJJ0XvpQ4nBl0zsdygtT7wTtFTHWJCX8TLmSxZtSwn68Dpp
7WSYBxXRkpl1LOb8qGR6c3OgfKGiUCTjX8qtAhdCbPG45/CzTlsHwSpHahlVp3OusPjgz5Hi483T
Si63A4Msmx74rcugLUhGa5bLCn0+WS6xXq34mXbMEFQx2/FuPhzgicNlcm7LSLcO/iznVzwOzsus
5EwA9eLyUOOAtqa9mUWBLtpwHKfM7Mvx4Ba4jrbpOErXDDrVuVWotNKke/i06TlLp7Y8MzhKt9a1
ygOB6EeWsv5qQaUPYwEKOrd72fG1GsIoDpnTUY/AfmIu6CgBq/RdMqJS7bY8rzH/RDc46Fzj451E
kj4uLJ6fiZPHL9NPwwDhoJM4l8N1e7JmrWe1LmgQDqpMRqCqOPzbocY7q4X5RnibjqrCa2ZnRXF/
6JY9Tt+bqkOs0CC2fq8L0E3v2tv1Ahq3O9PmsoLtf2a5uA2oksmN5SeMIeSQtLG9z0wCJnUIy9k9
tP2l6UvF1s/uXYFBtzPKhegohvexLUlZzOqMl2negH4ec1jY15szHTouVYDWw3enWJOuhf5V/1cR
3X4dY6o0sYPHUF5e0W3c/jdsAA+fdokjhq+W45d7X8GB59fngvl1EQcxfScZyM3UsFxMOkHwvTXq
FRFAir3VJmPO44VV/Uq31mjizZySQ/M+0c8VX+wJc3uGdWwhTtRdBQDvYUA8YG6nJDuADFmsqUJC
NHeXZK3GatwvictiGKHVXxKN9PxCs+s14ERGbkwzEKSuI+oBEHPMnDBcZrbTmc0i5jovqXdF0MLG
uppiaR4ALO2Ebx85shLEIpNFxsHgSq7rnKfVQG9d77kgrhAX2Ib3y9y2qFAl/usc8l1NiFOAOa7B
MFauWtl2tMYO0s+ol1bOEr2TbPH1b3V11wJXyg6kBi9CftLbfT+mmaMrElmGhXob92g3EcuB78US
7cwg/KmKfN2jLQysi34Jyu7IpaCvPRCz5JMTncElnOZ3IBg9UR+55e1bKlbkSe20qgjZ6bSGvoOV
E839Ze15u4t76IpoFetiEwbj4Tq+6pGI8s0DSouOhyWCN0BAe+kv1GxCeWN0XDAXEGwUJ70QzSIs
MDTP1w1+eO3T/eWjjoU9HxWD4AqCZXLOHHRBlTcrfKhBRvpJ7LWO/1GZIaZOJClV8sQAOOfSMDD8
VJpiWzolbaTVigam7sWsAnf//tG/6WFStNTZUEZ8d1hzMTQsGuEkEoddgHVbxgh+0FBe1JiXH9v6
HcUZdoX0/SqJWaGJS4wKwh3ySoG4nAjsqIagWZ49pjwkMswWlyi/77E2fjuQBv1x+KLt04VtyiBG
PobPzMXjdfAno1ycjbop8/ApTqPyKZ6tdUOigg4A48dR4aIgNl1NB/yt6G/qfhLqGbyM7sjl9YX0
MikCD8H8z2dfTm2GedxVyodpYqkNSWA28RDJv2RsssweQCN5RWR97a58XnrTZIGGToABQHo7ZCdY
s1pS0KMiX5JVNiAfZ6fEZZLwrzlrSUNuC9rnChCmOq1vwxn9EjQY27BbNQE8NrcxC12Nv9MRBhYi
t3vtuSd4usJex6fbVBZ36+wQdQs846ixV4FZEo26g7a5ZjsmKNIBfEAK0jTaTivWb3W7BcOw/uo2
c28/5Ywq9XiCU165F8rXD69VBhZizjlGK1C+P4q1E2SjPuhc+mgwzQZtOyOw37XhkonT3lK4Ikrk
6hvx3nuVojD1L/1/0jMbZKD/Zn4v22ZAEWv/f+L09ZSyIQsIGjH06ftoe4BQkJ4N1sse/lUv9Zfx
2Kgzv4yYTgq4bPM4lUoYpq5XwLmCQ5Ml/jHsu1miMIvb1BH4PtcD04mH1L1bOqgFQDIsrug/m0XA
csndWYl3C7nZGsHnnsLVR3md/RWTTo/53bfZs/jtEKt1mIsk7RXMDC3wPn8W/ZJfJ/W8ZhWT4mcT
MKcqXcCo3fhctXpmE3j8YyDwQZoHTEF9+pN/A9SRHoTTegRwqpFXe9kQTmUrZptOEzV1DJrn+4LU
27GUlCgb0hmLUxpuD9pNG3AiHVwV53wn3MyEwzDzJkE4zQ2iHCXsmzZh3je+aCp8aa1ZrVfQSsZC
rHsbVH1qqPWAaazpuXv6jJ1AKbRCKL6/qTowaioZD9o86hVLALkRhleyJRUpeQaGiqUW8rYN90Rm
eAVSKKVLk2fwy5w3VjuholioFux9JsVPA2FB6XQ4sLtns/DklCf7Z5Mvt9sd3bRhTqUji1OiCVd3
X0KxtqFZJfb8g0PTH9ETK3kFykquQoIVBMTOq4wG0bmXKobS/NS64bQTLXfChY25ZgZz+tiAWoLl
024ZiVRrqRXMn1wMHlcOJEPVtilJsL+1Y9WmAzFMqlXeqto7090+i9KLPbysf2LFeaVeCGyNS4bw
rZ/zgrlmCB6SwLNdgPbeXzObC+IoxsYQt5G7GDnwZTRuFaegdWKb3O45yq1dpAaoP2fVQtNB+bUC
rluNJsqbE78nSCgnL10/4/dtvI2Tz/Q/1N/J+CgRRIUBXol+47xFWNzbL8vx/4RZuM1pDx9Hkz5O
4ayllgaYsAZOUXvBVMrJyp1FVsCtWoGeYqZAICWGyFpQNwvlGHOw7gQzHUB/IfMuRHKlLsbBd8IZ
YvjoPAR6Bgr2/u46P13ZNGV+GsrauwVeyAADTJ8LGGiYXDQsy1rlF31Krj/6ywroNLOqvSVGPZDk
YhcJFI3kETgPqhmXU29DP1+nMZn1wiB/A/kPujd1HezeENPdXNygyhuRIhpD4iohQvEKvmUY8nck
XwG2as4JmkYY/rkcPDnaGkjFH+xF6v2GugRJG4aTKhZlWRvjHAYgK6ky5wt0JWOYMFSIyT6hEUdK
YIpj94aR0VlOXtzDXtTSSORhdTpg0ILi/7xBo8DSsaNeguipx0Y1g4Myp17ygfwHJjesfmmuRZ9L
52TNj/fubYUNGk3TtSvvWqaZK9XZU7HGMtjLL0oSPY8mmnlKfv6ZxMl93RXJwc7IUDSv/NthfZkf
vQrOtnWJ80n2F+nnflT9m+RN1HjKy2iBLzAgFdzsLFWSfrXOkzb+H5qgp8RBR4sAKerzG13wKf4F
KyI3aJ7l4w2Vlu6l+zss2cTPBp6mo4oGW6THYzTK14HcfWaI5+ZR0xeW6rMFLJ4JT7S2Blbo09H+
tEXcK/Fd0vWSFF36S5MU/Q4scvjCDYncq/CD6+fRE8RUtE6FE1ClmvxfDJOdb6BbpjF7RpxcQi1Y
Gs+M360BFMQfMgidwaipeJXY3E4+OTpEqRo7HfbEjzE3l+rZ9nFXbIZp8XEg0UhA8l/0d0LDayxd
+oOktNN+l0v1B7KVw9VJ2z4AAZWtQbMRGUxJYdxm7xtBxOEMmAZMPVFwGzEvvYzetyBnJE2MFR4Y
W1T4DmEqStR8LBtQ71iLvprsBLs8rkI/8fOdzL2Av33YA61hZbSMBcXjfxuiK+EwHukN5clhylqi
PTbZF17KgmJXlzhO3vkaIYq6AyHt80kfdxtr5B37li0uZ7+5lrMpmkM7hERiGoMpE57hFzecs/1y
M9dee6tnIIxIdHDMxQNeYllFkN59bplO6vwt1hwAlKIYnNTZS1yYxzK496yxM2N62cI3ERWiFp2V
L4gsxNIhiRfdWx54Lic6KWVktVUbjUnTd4Bst4nPmAvaRi2DQ0CgL5HMkCrdIwh1YkWHDBr+W2hc
s1/khHZGMoeu7Q4r9q1+wU4vj3o9TqTqZmkkp0UsxqXi4CxvwGuLgZ2i57nVVbwD1kq90a+9CxSH
y9Esyx9+XREMtDW97j4MCt7BU+vLuwb0HYKz4JGkaWGi3GdCQO5c2DnESAH5VYkSoyxOibBmjb8u
pEsUb2sSGRrckhRR73GFmyHFGU9J85QFQAa/uZGsSNiCG4dYUtozE0S9JuKDXgSyuIzbkMmo6P2K
AlICsixJmAdkFkaXQRngKW6cduOh4J3JJgWlWM1AyVVFt5csZVPxzw7BdtU6NVv95OPZOlDqjVfX
JW2d0vkl1Uoh7wfRA6Qibm9ytLuPYsozzzaL4vLV700FQI9iEgt/rtEuZqO9JVOzrBT9+ebPwzQV
u7WAvpSU2gyQ40yopjaC347QAAis3k6px7YViLmMO6KGZ2jOGcuWtrUxZHbVyWLecsYIJ2xXgQVf
t9fPfRHLbIwzpUfo6C/j/qkni3mD2OF9A7vya9Kk+CMxHCzKo+axrTRyl8/yjhodM5pg7rdUGHhq
XdmcbqgAgQ97mg9kpTXeI4JikXl0ekZSFmDmNk9emD5kIwpNsl4E3nE4kDybEiOlHAKFb7maawWs
UplXs/tR5Z7wzDlhnWI7bQBOOAgCF20cpcGPAkeksfh790D/u+ULFKSerkUpSIcZcejGYVeW+Kzx
U0n9GIDfg6FLxcgUvQLLw9WCZ0aQp+GjOJCJyG40PNLuBd3MhMJa8fN0A7sCST3bO99GE4nIrsZx
NMz5/0IQqcuuDFF+VB/J1f6levVN11Uqgq6h5kqda97EBiXgbR2fuN8t+kTt33hZVVlHtXK2vTqJ
sVYVF4hQC9kiUG1tRGtu7Q7i1jKY2TW68tSuJNEx1eprC0OoE8yOXuE1SqHk2Yd/1yQK40+cP65H
cvGIQjW9XdMAzaWi1iqOuIaODKR4lyvH04RScWy5G1JvbB93xqHOtL4I/EtCy8CCA2zPzcNAbd5V
sbEStcRVemnOK5Rdb2eJntn/kTlj8H0u6Rmt040qlTHyYnB24lcM0/x2hUIlYEnnyAcpVlj4/y+W
+nGSFoWNqhYm/oTnXp7giFz385uC01WvKHnVIXr9BW1llAenEoRKLEnhepsjncCyktNwMSYOr3dm
hnYWzEFYPC9wBRRHp+CvGzRkxFC9wnoumqo0nSOtBSZHfygVzaCH8nmtiQWDWCibr9lo6XFKO8iK
2EaM7Vz3AX0IgnEza48WkAxDLireq6U0bPD+v7fbioaUeVuEaG8Q5Hqwg+EseYBfEpB8u17eluBS
Xo5QhrFCAN1COMv2x2A5rvE4Azdf2jUE6JlOzOOicvSEEWYWB2wnHhb+ujOcGu7qHGr9VhicGTd9
EcCegoRY8Igr5ZCyHIA5Kkaxq/EQuJxkp8ts5OzRqOk39EAlkMWE6l2cm1kuj9MXLJvWGt0LkBZh
McLQF2hnxPCfPKVIEy7jgF0evVEM1pKKFowShlbmbxwrk/09Zd66XuNHw04ooY9TmM9fEsnUYGnQ
vCJugx4JZ7IZHIo2xS/0M3qgijWZH9m5V3cBFCcY2QvfLYhmgLe2gQ8opoawQ7VO+TPG0PW81eBg
UKgUfPctVJoCJJxlGbsAEpVm4t7HSgm+5A+kBhZSG6YzXrJx9B+dKu2YpxY9CChSSxnWntQzrSbO
KVX44FSgVyDHltR8U5xsrU6W/A7jwf1CyuTno9mSPfHAb1fWRhzbRHiGdye1TiVeWYCaV19DHkE0
NGnx4Gymxk+IKL7peXPxu8aVPILUIMxGA7NN+t5abegQzyT+f3rIxZ0yUamepn76Y1twF3T29rrJ
novIvdX2HXANrVyPX8nEhiqxvDekHfuW9UcgcoIqvRYnBNlfyZjeiY4QNsOl7ZsYNNOccSPIRNW6
x4y8SrLsv/bLUsjt1TpMByWyee/bJXqbSzUxTzmiz+29CMG2RQ8fj0r8YlIdErDw+abrgFldPvXl
9PJMkfjSAieN8Kzp/BMr/EY+N3fMXlhYw+1W57mLsQ9bBfLmS+4MGIhWXEWL5ONAKXgSVdDoSvo8
sN3QMdgKw7QwVJ1ZVZg869psYo+Q4DuKjvle2+NHS3QB0j9+FjMYFpO+yqhVQgE4AOF9ObizbwnZ
tLbt2Trhh3YYXbh0wjFh5CGt3NDbasb1iVR1wRnXDtJ8UlD2FpvNQmJrfwtJEhUV5T9Qf0CkD9D6
CQF6Fs5ug3NLaLBeAXDiKbceUSATgtXTgJOIZRTReSvT5yIypEzHiV8iYkh5rBgM+mBhTA1rb3xR
5V38tNNJiwIDXPz43xNemcXy4/82nEeYHP8oPzt3mtdy9sY7lIKvaQ7YUXsDnxgRr4m6C7tA1Q5F
7Ns/3w4UAB4NBCvFZfi1EwnbwtlLuQINvBQjwsVjMzlRoW1z+WSxilpw+k8D0+Hh/cVWbD7p4hBL
dL/QGL4nuPgnT0IFZWXJ/4czoDmxwq1r4fDGWnKdxvG7pI8qGxfa+TsPOzMBKMUyloQM7c6Ftzq+
ll617zxjc7EV4ckY0AQAf2lCknDHGTrfOXdl8SRoxjL/+v9iuX5EY8Tr2MTy6IbVVtW1LhV7EFsV
WfrfrB4CETb94d3HYRevKR7aAuFGDWNeIfTKdunrKwMLJhqk9ALBZE6oWtEJXMJYayvPgJE/FHvD
9WYhMWU86KnWRJbpzwe1ASjhAkAnMxnro+gDO6pWYAoI8dzTsgJUpR3OZ+EcSaigffbh4GV6bPxa
H5hyD+462jUvzgtMkrqrlYWfV0YO3SESRnOCELEJeeWAWojU80M7WgHfhbXgI8I9Talj4pn8xnoj
UmfpSmuIFY5Hj5rMJWPbUUmXxXoYff2kcllyJY7tFBinY/WgZybf7DyPmS8Ki5Cc8l40YGqwxTeU
fy+QIwY49m6Vdx/jwp/JJ800qFbErbmHm2pKSt5jsE8CnXzn/zTp3edcd4qMbWd+DBoHff+83fUG
8ISoij1ID5B9As9RDlZOrVwEx/Rtv8EUp78wQyBjq9YnIunHnZ/y71C6JNBtHa/iWHC0Vq2Y9Brb
WmMkVQVvzHLRSxuZ1gVIO7PVYiJRlaV/lykbREnbo2OEiOpLl95n+YAlUnO/2glq1g1RyaMlkqMO
dza1WCgFefv67y6S+Shw9dRGdtMJWPDf9A49TlI3EfEc8TIaMhPUbxvTJ/uQXClSW/uz1vurrOGK
NfoDwCk5e4FRUUK6OtbNdyc/ChCGwsyncoX+pJ952xoaelLViZ56CwX9DahzRd/98Q9eV1puLgQO
CTEMVKr5NavqzMmPvIth5IY45sm6FKKSVXPFe+0N5JUZ49A/4cFC0w/uL6+j051WK5L4ndPBY326
ON1euxGlnc+TG01yJec6atYKCVFhFvR7/3p+HFFlcP05jOKf1MKceCi182ZmCUVgzPw6RX2IBje0
tsoGp+08UjgKS+QUhcyoFq6FNNK7zsoHm7bDsMS57xG41iS0eTnPEgMi5zYEUEp4qkCctzj2746B
ZeCKu46rZyvGyc1jY06fZEblWTpJM0hFy+pEhMdB2R5Ib0/Zf5QrN5lc+siX1PhqXyWy8DW9j8E/
Ke/chZiuri93PiQlezqMPP3OU6wKgGeLooVG0PISaOSJVefPRoTC65qtfEJsvA0XMJNBLqst4o/I
xiGsgygdiCFzj696xlqon76GFnTfvZXbqKKxzwuNDqtPh+UTZe3SME1T2DK9sM9otu2KheKG4Sdy
I7po+cEfrmJRbRNOzGneISTdMEoEdFJJ7uzKMDsr1Tr7AXDMAA10da0zejv5ioITzvg45/wc0+fw
/g26U5/r4igF1pYhgSMsMDkBL1WLpDWxGSd/pUFqRRHmdSiAA6ZHaMtAzMqkVy0r3/X0/L8NNN6L
W32cEZnzcEviZJszLgKC7b9fHu4Tnfgv+BqUcwh5lsimxXaFtW33Z7jcH48xHNxizjFNboortdLJ
mEJZKFv7qK8p/Rl8FW7JYB8jvH+roNqdz96jDFIBpMO7IJVdDWRPm6Qal3vMSqoNoDGRwECwdBG2
rwr2rATjA4cywCrw9Ubl+NMnIqNF25MWji+ueCpvujKQRql3VFLcp1R7c6UsCzS1Gv7t6SKb06xO
7mIMaGKIPgKNChs9fyv1YvC5QP/H8LOCtgYncFCA7AvRyfPstZ3OUpvMiyC/mDuW+ArZ8uLpqKZ4
arDYZ3TKi3QgwybPP3nVqwjdz2FTRZ8xAIrrg6plIyn7ddWiM+2o9AIOguV9b9xZow3hzHqck/Ir
3a6MuCuxc533KDotGuso5aXRXF0n6Zu2LK5ony7ddP094M4PA44OTQGXt0VHugvvcxS7PJgzpBro
9qqGvC6qxgY64KUK6X8e5anMwu/RNjF5AI09mRf1gpRzuDKOcLGhDAVkO7dC3Tw4ydBUdmQs/95s
Vik7PxuWMqhAREhKduffthJ846j5z0EumWNC0m31Cfa5Slr6KtubrRxlydEHF6Lszp5MaoHhTo/N
yeqK9vb8ljgm9eNd4vrvWvDBZSoN/oGF9OU/N46l8QNpdqRcKZ1k7kn7jpD1JIP60glDk3Kt3x0C
J+ry1QJNeqrpKYXdEXnQ0OBTB83QN1VAXiKI3Opyuu2ZWS0Nskp9AdOkVKbfzPUqxPWtV7vJWYns
2iJ+YIscySdQ3TMNFuJnyEeMt0cYY44c+xzalHtCdhvC5Tksxcq9OR6AkxTLCPZuvKk5dDzyHOTP
VTRByAO18O/6WPZqeir+7eJVLxAXZDfMOh0HtJCF32O1zWU9LL0HrI9dL4/rCkeCnv45w3qujrLB
BxRKu5ece2seNsY6VZ5x745WbSYUk1jNT6+dUHQoEhah9km2Vqi1BqEIdDz4VXQ7CYDBxExPfdSi
9wXQ8W2LEBabmZt/ChE/wj0gw1ywT6h7gtDFLab183qO7yXHeThPLANeexCuavOMKMbXXTkzjdA4
BcmZWNlnFgZwjd16+4VKYniRJ+xGG/RPhBw03USqt+9vZggY7hufR/7Sf80N43nSWtpNSqolCDGH
iTW2HVAm9bkmQLjJt+RsFQQfBvlvr3j9kGmODZaHSc3TvwBmG+MTlV5N1O4N1ea/Fjti/RBqTf3Q
zED/zOsJS9/Pz+vaOKh7Y9/2nPi2wvQ9EIFh8eE05nFd1/6W7dSvIwJVeL2TBZ1QXGgTCOBnd81T
ejmg5diImEOqISKw0fSG7RuHr6/NuAcUioRhR4iCGJEKlNlKK07ddJImVVfXRje8oMLta4WRQvvE
WGJpk7mF/d+/xXtWCazIIJ9b8H1Opanulf3jGiprLpE1jisz1Kj6P1vFKa8uoVuHXWiQQmtZYxhh
9k3TIX3bjbdQmLv/JS2TksocvpJ9n1qbWGdB2RJS6tU/uYftcal6DtsTl4kx+8KwTFzMumhpEcTT
k+7ePDixoZ05E4kICbneV4CF780XlEbsqKY9hvRbbMUSycjmV3di0bqwL6Zbr+3OvIIIfp2uBnE4
uwusxDxQSFMMjWthXVDV7NYKYqwny3PC6LHMM6FLVO47sMFRwHhu7OgZY+4MVLPwbK5ABlvjYcko
nzGq7Vu92WETowAfVCXwHFLW6Cp0CFSpkXIeRRaBrrh+L3h/lFOaoSw/GIgM6JGZyyrq0UctJ7iG
uqXTKRWs9IEko4JpMBXhgmeVVT+8K1knNdHNT4/uTO4Q/GomrfAPxmB6JPa895hlpQoDtyTClGsT
lnfYSF+EnMbS3X9MCwEIKQfJifhzv84NNeT0mli7etGbWGz3tt05I5dx+1P92xahxjpfBBPG6agF
EJcmPfWdkZHBQM38ZmvQ/R4JTNjCv1psWi9Dsb+quSuaOW9wQwZWCx8xdbRFSHPuO12DSR+m2vrh
TrVoRHzp8S2GGtmisK6M4WyRmQcJuKWSQ5znaPNj8YxsCqRp6pcARqg9KZv90OF3S9ZBYRhzryvA
6vCh/2dyq8WvkC+a+qwlM7N/8+2gPMEfXvGTe/dSMzPXOc9RCI3lCRsyYujAS15anOSdouniJPfS
9J3qzMqqilZerQRbG4sDX+LrITuytw6+Yx3G8nVlMg5pumcbFH0koUeR56LutCzlVQsZ41Zo5tRs
WwFlXHvp9d9zFI/8hI+4cahiFSl8kHEGhW7EdwJ5qtN7eEkOZylIATuBBsOJYHPrrGRY/VPZSa7m
RKZxqxRQ5tCBNujSP2ayEb3qo+5Sp3Ehoe2Yma/5J2nkFY07NVV4h4P7+++BQ3yZrzdgQj+CuBPM
luhka9vr3LqmC9KXgUYaqV3r5TfoFDcnNLeccQdETSYD7jUpYnEMnheNm0A6C2wbq9ht9ebeghwu
haEO4LrOe1Vc4uvNKduRke7VOoJdxYB6k4n+9YTUxB8se6pr2yY8RBLYMarHBiiB0saPvBRGK+/G
PhkhOOzM2AlTGwtNl/iXowMBrd6vFVemSHzm+jIv0T7mOHSr+fDGIud73uqrJJ3GsHmlMZaIefx+
QH9zv8QTrK0HSknzNv6MPmorrrHg3DKG00BDV91+iigRiL5hEhndH3GHt9rBrBe0bxoya/IN3Ui1
EBggpcEVhbwfugYK8QL2x0fuPXuUhuVNWWp8Ia7Ytodc/MJAWVgGjUHt7ig+bqhsO9NMNhep4vX6
/rk8n/I2kigs28N2hZPld6VR745QSBiYHKwGMA1Zwciz06HMI5KnNMiifED/pgq+WKB2OZ6R4Aff
82wizJ9flTLlOHRKZVNQX4j/I16m3hny1/MkwR4rDySHMTMHKRasOk13azcri2y+dM+dRuTVFwCH
8h9zcWuoOXWW6RMq4cRid+zOa4KUn6Hx9WvDzoWYkIOcqJDXCq69GJmnpDIzRUka38N+5yQ7aGUA
7SHsxpWuAviihZ1Hxveo1dHBtfLOwgpFATCYl68XW8hIk8tFDXYAxx6qxixOqByH9soNfuFeumw4
vw93LbPcUnQURoqFWwx0JvugjXhcLU0MwhvX0S4DN2sGNbOYIyYmGCnLm9I/vMuu/bMbgVnQ+X9y
XWcc10ApiGgjLV7DT6EIgY4w+037pHfxH+cwMu7VZA7Svhgretl98j4W/MFwT/QaCKDM0ewYxlsD
MljNeg09jthKrY09VdLx1Bb0SzXeqIs7mU1Pk/ncSgVVPTvh7O9z+3MZuXleWtYWQzMqA9ESpGkt
B71G9o4YIvB+7319xy0wwKRUANrbeV1jU0JPdl87QKui+SnwvZpFjFU1ZM2Z5pcrIiGezK9EXr6B
p9gvb4l9CHp7tprpw8mpT+4Vw5bb4dHdkccGrmyUuYjrakUrdE22I6Fj05lojohv9i8xcVRvGO1o
Rub9Piisin884OxkJA4LrB4lqtr4ivaiwIuHBC0rXpNE+/wvLJtar/xxhw3xpi7vXrNSE5mPs4TQ
tAUCmffOew6MyL8vNbE3afuxkOIS05PLM8xpvilozy+azMt5OzdbEh8sUmAkB7vnKOs6sRYSvBQ9
R5251qwsy5KZnYlT3A3mrIyVsWYOg3uw6ECOqX80RrRpPC/N46nI5hANW9C2e46gjSkC3Tw9xJ0F
clzCtCmMNGDYjzDgjbvpEUUWpBQrgUFHCjmHpZXDWQLaXxaZ8MzsWBcnXSAxJ0t67LMHeaLgJeW1
CbSldDZLihr2hqqlHYEGCNnsuOhe7Y/EKd6Y+9VpvL/NE0wd0AGxDoIixlsQXn2CZIVCDrDa1CTC
hFaq0fogEThe+++saETm8VdZzMsbRDpnc7HbFhia+woCz5AY601l0Xn8yuMnChKpmA6BN9499UV2
4ePx6HmcQEuiSQpS6wQPQLnnKMfejhxalHYrz4riXPmBwLVnqfNYX1kdWEISGpb0i+nnJiONmxr5
vBEn6LLtxDMuEa+y2GZ5lpvF5tEWzuTkQgR3opOBtko0QsB4BfMyVoUTUU0k9gXn1F8aXRXb6CdM
QM18AXdG0L1lrQ+rhuqmQlkG/8ek+g8Qvs2D+olMiC1oAXIVYQLNyITTYzSiGzFo4Q6uj1Gh1iDP
bltWQfvnOsO6iy7QARieGHU8xt+8lJdBNmjp4q7gJFdH+xtPW0dqrkmi4xm9Rk46WE8bOrUyb3PH
o9XWjyAlGJs7yHRvSq6jgxFU2gd9A9sQRTKcGHD5ygRXQtBpJfjZWmaxdw4TCa38ja/Lh5GmRMyT
dE57A2oJkgwtMUv5wKQjtxG/2NgkwZV5bwsGP5gV59rHuejbY+AmIGDpOmErOCUQeC+qV4fDYflm
Bq8JdyPbyc06DLYjekjW9S7z2OxREawuv7OeQ99w6uV9u3ZfJx09BqCBLv6KDZsyGnb9yHI2gRKg
4ZRvU/uKRlhdYFdw2P8rXp4MjgOSKRUt/+VCCv9l5XH8cwMhJEwKTCFlbsG6Crz7fTrZW1Z7E1Dq
zfJ+bo1lJoEVaxNTJN8DeTcvKfneliSGSWBDY9nQovVTMGl72Q1RATK5PU6xQ2taQfGSKFIS0lvt
Mbx69K461kpT5NHJnU1ADTt9nhkCaNDMND4XiE3bLw8KxEZE+iy2GwGRNx+bmfdrtQf/05kfdkcn
qfDKeh39E0AJCD+Gp+jun1InUoJ6F54ziRR1zb+17YtBCM4MV9h1S2UoGyLi4c8YDUXVijJhGe0K
FH1i2cJkWGtzNynk3BscEXt9PCbYHHsPU3zGAD8jFWxQ5M1UxoWz0F8S9lDO5UofeUa3YYzWWSpt
nrDshaDNm9KGJ5Z7UyuJaOVXYqK5Cv8WcCnJBbLTwIpreGZFi7uP3CQ+CymOQRj1J64COk73ZM2D
g0WC2kDETT80Ip+XWySBToroM6J0mkJgWSf7dFnASbkiZB9bjZqOZTL3IpFhe9ibig646JZvUoeJ
uBLBwbLRBdNxDlNvka+SgbaWhBr164yOHqTZC5IFDHqEJIIo2OAW8B01sZUhy9WxaCQUHorAUHt4
wkM9tQmc+PyXhSPC9+S6jTjA36TqKUmcEzgd2CaglPXIK9xtZpg/lsUM3rmxlTfxVe9XH93j/dvc
WN/GJHGfyp/i5mdv2p+M6PdGzq2NKfl2no+tObUXzVaArr1Hw4WeuZPKbyZmJp4gMnInkx7wBLf2
THkBEnOwReYGAVXDcuOzXAcGMH+zt3HwSPKvR4aKls5l+dPtTJtzeDS2UJjxPVrHzF7uuxGoYCWc
YlCG8LPT7YoRAoYKQSKF93YzGhO/KIiYYLZQuyOoZ6ieU33rOsqcPpHMA8T0ICA0IQBwxC6sfqQX
qd5WQnItKDurrLg/MVExUKl+bVMCw3V9aO6G668opG3slZb1HdVnFnek0V4U6KMC1GSSkqQcppBg
EYH+omZDG0a+cAdwF9OwpNhE10ufyiRZoNvFon1D0kFhcEgZ4CsEdB95mKw2adT0BMGKXef636ZE
ubLjBk3UPSOsFTH5pTC8lwne7JtEf36ONEm/hgTA5CQN485igIbyPe2yFmsZj5wu/PEKb1B/nCSS
Ia9sbZIFfx0WjpPqZxrO4zPR9gWjwCXH8ghymkDIzm1jR4MbtrBUlRitoaXolrAoBESJODkxIvWe
E7kY4IlVl5cwsc0G7Z6BEIPWTFMbkRYAih8bHMQjtmpGHthFTgqpFLHQdKtcKQgcVck5aNpfN6lc
TBvls+g1+i+SESWFhV+khXU5TlEPWochG04zfrakoVP3aOpcUd3EXtjTblkhuo5a2hdzPtKd6QA8
jcq9jiJTQ/buazRs+BMb5HycD2Hi9XSzprsXH+sXuJMadZXOtAe7EILg6/BgBQ6xceWEGCAbrbsd
06wkXdWbK8+To1zlHBmPctFiqNfEd5alRBrDt7HqxMiScRU2IpRYkKurGtxPJxD2wQwFlVKf851Z
/GW6kb2r6+2bYS7ugLyq/Zn8o2rKPXR1o5HUPooX4N2jGZBHkkJlokWeRlZHCIpKrW+Lm01ZmHY/
0dfG0UAAwoIGVue6NaQHnIKRFmcRff7q3GmH/Qc38/u/9dIRNUO9ZZ3J5iahCxSB1ZwnLqrGdJFL
P92bjb4Qyxocbz45NcGYulERLdpC3qeTL4lLP98XlWHTthaIn/6KUS1W9evW7xYQjBAjxw3ikxst
jpAtbeDy4xxbGtfVzWC8K3mtEiWJbMr2S8VmSPOGjpb/h4+1NSswVQuo8gCH2aRWrMH97pVTNSuZ
0GqEkD9iC7FZrBXaFIfSujos+3xDGbf/NyUhLA8P7/p11y8E+4x4rq39MmeNck3BSw/rdQaslwQz
JbX7NFWYlHxLaL3c0V6qj76znmaMAjym7/uGmrFHI65hEX5do41iU5S0jGYWXgqOy508v1QLvXJL
7P83tPSSOM9CyJgu97Fl71jmQ4FSqGwwWPF8+UhXwlLI7LDJEtUXdU2svpkyqZ7tQHWQ1DWL8/mY
mxFk7MJxR1mDrfVAxiOBaYzRe7hm3N7kvJ2I/yTw4nEHQle4EA3NW0YgnYjU+v6FLGfJkXr7l5SQ
PAtny2FO7dsRa9cogGorwBzmlcNiQUquLulQ0O6Osa+AZWlugswd20022YgIz/nOREgTZZ6ljYig
1vCdyubH5eOlHSYt3i2wd/FIAh3YdWkdhFNfQ4lfjGslAGD4E1eu4Ss0Nbccu0wn/XgTECFQwl5k
AoQ+1s6xTXThlGQiP0uuuBXuZSIzTZo3UgoObrPU0/HVlU27zqJzxUd3Zb7IhGr2eu7T89qLIShZ
mfhtOfVf8h+jjXQNaoq3nZkLvkUpo6mqO68deCKsEu3C6Q+4CcHlgoykmehQwOsRJHKyqImIW5ka
MgIyIXxx/4OOq2U57ti+9wpd3nOnzFFKxOF+3bihh2EsuANKlUF5uTr/ywDZZqw7sKA0nOdJSjNI
qKsTp0gW9UmxULnjyM4qge60abyaV14QTwrLKd3410zEX2xDsOsrZ2Oe25E8aG4LF1ZvtX3B8FSa
UvDwHAux687sbraAjCTIOtqdlXM9ZUmO8v6ylBq5PA0OG9eFKe589bQiw3KCoumN2GFQtcUi655B
tQGMwnqLZFTJSp8T3cGkUJcGk3v0fRsp4tkVRoOQbkturEDEHXXvO/RIhLCi25IR/E2aD/Ml7Bsu
IrMQ4r59Nd82XXy3wL/Kb4JPhvKvadfEBfaH7OampMkAJIByORUDFml9JvGIewbbhrfZg9AjVlbN
TKj8Qb15SzXzPaAdtbkcMSW9IfUAKpEO3jLaKpXMoYTptYOwCxp9aCXsmFOzMMsK6aHb7trAj/VB
ka5AdeZToANwRpbrVT6/WtlKmtflKulJYSQMxFKZJktn+AA2/Ba+3Bn/4LzGiRTdOGq/UttUx6Rc
6O/TfA67yFq4v0jDiJUcC2ausX5FISCUU/lBzk56h9R9ATmajezDSCdP6g9WJWeQFdMVgdBsY9Us
JkqF8wX9arC043F3TcTctebG9nKeJ2mXMM71xFIe2r6ANZBwhjowFHQuDPS+8x6A+G5t9Xn7Folv
d0l6yp072Mp9ABvDBBga6ZEhnpne44EED7USX1KQjDasfuoC6zC1U4f2OElpOsPXKgsd3nZMSUQf
MgD3DeGQwGEV/ij4hyOsEN/jyw1/lhrDPdR6X7m+kzboXvFR2U2s9sK6DaUPYhGKPvAz5CEiZI3T
1/26DUF9pcuJMU0BAbXkTaKDXULfkjMSynvvFQi7GVIvxkg++L/7grFkS0aLWeSvtle8P+uP45Jx
JD2/W/R1+YJwrtJupYF3YPYPmSMIHpDQyQKi1LZBOCI/bK3gyRwrT997Lc+x1ogIpKfAhJKNQs3c
je6HiH/KwR6Bwg8Uv6z1758f0ecdyuqrms2PuQ/87HKM2n1iJ45EXorIsZTqOZAQnLSHWwZqEf7b
wPxwRKLYVMV+3FTyJQgauoPMYhLLEJezuujhQEczz9kwiAxzV6DcrqOdjrovtdWQShYIHgYSYnbb
ZjcD6vMwjDzm/jmeDlhXhRkWGdgMNINkeljWorlNzkPKPBq1+vfO45NZUo7/48q6SxofMTbzt41z
Kc1mYzSgxrHq6XdJQsZvH2eg9SfDmzhqeVJEYCkU/4vwlP7vH5DW5udjqwmVNQuw2PlhHX3Hdojv
WOzThF0P5WEiP2ylvFYnnChkR4I6JwQD3CkVbk6ULtVXYIdEi6pRQmmMVjmMLNRclFhmkypUsmiS
YDGNBtGqi6J2octejsmQh5mvQJmIxyhUonORM8c6s6vrgz7oFxYZSGDWnk6VMXcu6t+ss8zWLOTh
GGMrxZo4oVEWKpLpO5stBSCYejHOQZ2cQPcJ2CWyQM5YqPSQTYe9nCgVgzU6T9N6K0Jhm4bzk73p
gHBf6YMYGNNKDVhB+73FLXublQ2e1NqrR2h61XAU1LkYiCY/L24MK2XAdBlhadp4AKwy30+OoAM1
zn3hl9LPrby/ADcnDPR1YAaperw+dziL+aoYcAtbe0tR8gqgfjts0GKX9+z//cU0XDb2yPX/c+DX
959Wd+RcmaoZNEpn8WhxU/2gxFN+4Sfp2jhV9sLmdYtB7TLe5cZvqJWDqMpwagiB9yLNzn3DMiYK
hdrV7DR1nykh30rjws8HpFsivxD4EfRW28qMH4UJNQO+rgNUIqZvDesImwM4E2hNUCxQJseJ6qyA
uY/dwTJ0i6H3ysAlj0bXfKskppIqMTj9D4i1JFURJiR798p9jk3GVl2+Gr/NyfjSqN/9seCRPnFF
IHqqMrNct9aMioNL5tvHWRUvIkVwiig1z3C9JPdauBn7ZnzvzycB7n4dfZlbOZoLfk4HnBHoh9DQ
C1j20yIHwztREjahrDsYkJ5PFFHpzFEC6ejl72t5DxGz1N7sglpxOd2fZTQinwG/5DN13NxwLev5
POJf7FATSW3LfbqaHw4l1VOSdhuEkL4akzwmbv70P+2qwtcIibSikrKlPcwgYqmBxfqSgtdZ/ql7
UOu8uzxssghR2PoQ6ABJM4BRHtzF4Bn1bbmhS6X70NKFVweSM3G5gb9fM71lhWwcTAPcVa29uNBM
9+xgt0iIUiMmoQdyUl63XNhH8BBkdLOXsw7HsaZPeOgUVi7idJlL0nQksEBKTHqvhci056hzDCuG
YiURV9HSwlGlMgBd9yhya2HGiNlG8VjVvX67pb/wWESFNTD74Qp6hz6hIKc8BjVen1++DbXs7urj
VhkllOKFdGhL4We3H1SO1WlTmxnhgLqaX026wXXa10MCP0DdKF40KZSWfVp96fd1aaSDMYDAxOTT
vl7siKtlnzDa/kR9CXtKXnsJl6DAN+eCehY/BEQENOM4nLZcHMzR9AC2cYZnxGeib+0yWLUtVn0i
Gf6FC9wYTECv4uUYhPHyyQqcxO9rdI0K4w8phrrB8AcHW4t83xqqeNnIqjBi6hvggN8aeKKAeMPG
UPXtNuBG+9wNNC9UXooRjiFICKWO1+DEO8ctobx89D+kX0yIcY6kAQKp+VNWHy9PDPuVZZ/9T+Br
25cokMvApWpVkeUzoDwwWIuSfs8QOS1tqupZuZbLzbrfT3i7DOOguZK46PcJd5R4y8kNIXgT2aDp
fOQyxLokVa4mGUTrqfYWcJVxLqk7SC8kOie3da5MKQdDqLAVC8yFNiWPDvoTLAQcU6JDfWvTMaXd
ynirFcG8/MXvYn0tnuvBgig/kBW1GiSoAccTUxQR+7v/taEFG5/rmlgyeG4pDPVcU2XsaRiYFCup
hKOCfnpZ+t5HqySn42Rdw1nquLaozyqktxSqzhv5PlAFEsCz5iIeJT3iveHuni67zZG+EHPOTFCS
vZL0Cntl06H7Mu2Wu8XFWqcxsgp1mFErcvtuzjWke7vqG0j5SOfxzP8Pk2uvlrEGB6zJaIt07VTw
zj4V0xOU6TPL5nZ2eBeCYOgASizEGVa25sPPAmp0F48dcmI+9TSfCH8BnMZ6mnbAzii1si0obB6A
UR678uN1CascZzdSZ1sanxZNEtUeRW7si0PLJ+i35ScKVUsIcb8XaMM4kWHtXXZ5fPSKHZLx4V5S
X9LE6zp9U/el+tMJQd8e6zvFe1Gr3SPVNyeVlP9JTc7Pr6FcvQ4X6KfIFRlK7xzV0nOeigz8qcPd
Wwbkekezd4l42mR0bFoJCdINZkcZvetlM+U6Ow5Vc4JQXXbo+6Wk3enly3ke5EV2A4yRPttYVQKj
vhGCaCsREiirXoGq8PoK7+OmU8IXHjL3tAknoQa3cEhEvZV6XFG4umMhPdbBuz436rPidoCtyhVg
48IcaWojMue7B5T88S4OqPPiZzLb1Qatjsdl33f0BYWDODtU3zwcrGWclGNYCniB0KczPraXBokQ
4TuzuFII2YgeB+lt6BRIXlKiLssT+5ZFohZ3jEC7/4YhDKxdCJBBPV+dK6G8EaV60LhCpf8k0a6g
15SpvT4AJKrKMl3W0b9THRhS+tZzea8oofEAbM0bofHoad0WKrwTOcLk0lnkHLfaQeS2/JBp/v3e
ebj28Sl6tiTHoDm2RWP0DaeVC9ysRvjZ90x+dsDMN6TT9ORKjIQYUHzsKJ0ScFVmgU/9tqiZzMxq
UV8kRmTCnuxxhEpPpZEFq5c5Jvb1kKglUiM3JIEwj6EiFhOStggDj5yqp3sgfksm/5vsgXky0dGa
g63Xqkv/hOUpAB2TpbCpHnDrh/TJT3wrX58OCxTArxeIBmCm/aQGiY4Ydu6GXZh/pb40rzLSVNX8
fCLS2gRpDfq+SoC5TBoqhzykKX36J5TEgyoKaCb7qeJ+WC9BINEOzkIv23JswXcPM6WmElbg87s1
+fykxLbMKEEiZL9y8RZZzv3hFXQekqvXdJ7zCQSMvonVJXOJfPvnwAbxQT0cfN093n3kxOpWCDT1
8Mtml6zBbP4f1Jrjn1m8vF+VAX1bOANtMprTLBcDtR1w9eXum6IaXfF6EK1tGjzy9Y0mW+sqgAwy
5Rim4A9NqxGAbUVPJnmbgbmWmxFenbDPpv6tPDKwP8s0DD0r8tRd2fXs9eXRqXI90hZA/6toloOX
W6nlKXdn51saDsK1hPiHNsbrTayuw5uELJQnERH6hofWo38XNjawQIGmlndzX7N2ku11hZr/OgDD
Bg+0FECrpxTna9YPsXwff/8234VG5Hly6Ru5L9y1e6YawafATNPaYKoyCk5i9M/fAvWOMn1RysmP
cuUGTmq9JJvTEEqOM1ZreXzn+/i6bQsWP0j+JMwB/TVrTFmU6XFg3ysi+TPA23Y2ElwntJrAsOik
bgSo69TjcYoAKLI3ZUxjF9Mrx58lfcsDeXNf26nkvl1r8MbOoX1V6+pGaY6QLuA1T5VAD6O45p1y
vqiH0786oqB7Sm5cBmPQRx7bBgTvSAnWvU6TIo3eqNrc6AIcSiTKoBaOXM+pE0ONUQKE7sOntIfW
m56+fFflYBOJ5wOiLRi+7qEmHRZ1LxkJ3hQdCwQh3ui1EY6HMoG8+9tGNaeeMGldUPzYOSpY3ou9
M1pFWLtN9M7+5v9ARdE41QVB0bqctsXcaT8vu3bH1FXwv4biDRqGQsJ6FRoxNWDzzK/0h25QAxr2
V3qXvv6xOOo9cE9JiITHitbnMPL2ZzuYH1yksm4/+fJJe/cS59kjrjnsr9C1VH1uDM7T5QfQ1GzB
1LaNZDWWQbSjolPfyX4aIkUG3b+dd0UYtxOppQnGXg4gDSfg/EzVak4HWRYFjwovo4PejGpnKeRW
z+OiZhYIpBw3+WDdXFmvcnrf4/R3+HlMzROoeaN+ACA1mGIrXydHQQjAPrCuffeA8Ef/BmJKejfL
2ir+2Upc8rJSba0wXkLMcNwTyfzErFkkb9Do+TjNk/OL3EbbyvI6DSR2N3T8UmpdPmKzT8g3RiIS
+41iuNU19bMp8c4HUNGlPpl2qOd1dwtm9WPOlkENtMO/9icYksOKXZ6uKGgw4DAa5/Fa9xxktpoT
NWCGVDrkUNp7M8qmTqheKMjV/1CiNBPzsJSWYrwzqock8yjCZDDT0BqGbTSHHU7t4hwsCRarRZwY
vGPV+Y+Pq2NdTzWWFzZz3WwChs5UfFH2S7FUWOLTOkYZjE3ZVF13uYoPpnp0os4C3Pt1rFUDQ0zY
TpOtl/mk3qNbiRcRCkOUjQyPHM2BjviYN+BLAq1l62pUJ/iOgDBJVbmsBsNoAsaqooxsfuYm8SjY
BviwvrZeY3ImrjbrgAhpGgcLlqMMO/pYGLm6c2BxXRR7gyFjSu2XzPX0+JBo34nfpUAHMDcDFSAL
HS5jNcrz92nHwcbhtpU9vqSqWEXCe/M295VkLzIfGtwoVGq4np3mQy+jq7o8BZ8y7zlImEhgEKyI
c+K9UHcFOjeYHHDNIBFBoivZF6MYr22lDMVFXO64eo5sePMhVh8ZoJTQksOI4wZU+5Pbr7aFqCXl
/WflG5hfQyimH4nP+Lzzehm4UPCRUuc5ruNgQKdz7yqRw0n5iwbpxd5fQn03JSObkByUm7C1lPcN
eC5Nk3z2evD9Y/nhDBJuP2/T+cfs2ypLsNEY5XjNgkJTv+pOlocDD470ogS0YcxTiRnNyenhU8kI
O9WCj/b3BF4MA9rgqOGqGMTJIR0ef/wKrYaIKono22ejKOraAmA2IC9gjwHbHP5l7iouKIIUzPXZ
BPLe/ZquYsyM/ewEqN9dtinFI+vrdE38sl5DDlqJJ2NZu/VW+6hr3HL3CXBMjQBBkrWVjiqw6xDO
1ZoJ5IG4mtWfVoI3Mi3n0QC1OD1/CuTLmkeePBHTQTyGJMqOQIp6qkCb9z4zLuaa6vDV1H0gG/PR
9HiDjfLOTYI/Wwh5Y2hGT2b80BuoFF+ZTuU6vDdVD9ox5PLUIimVWYbZvbp6+o/6Sz4xlBNY+7ry
lWA19vjenMLr79kSF/GaFOSFFhf0QFSnQwILZiyGmZBkCGwESXeCg/xEuR7mcfLggrGiIeNkxkn3
6zDgIpr3fPb7vqA4ekkzX1J4h8nkAhHOjSAL7XVZv6Y4KChpFtWcn4kQ9V/jdxnRQxhzUsAG3EKE
UXTSHAq9P2T6umoNhIFhfFjSodsMSj6f2TUn+kvfPhusIB4JI3Gt+UuOyF9km0tAwEUbrmsLy6Xt
p5d9OMwuzcQV24A9OsYK5sFXlvsnr0yR2LFLoRiYelxV2YA6kiUZCZ23UF83YBYnH+3wZosZLbGf
YXp8sXTIpYFKQ+o+LCauf6MChwoMz98bYtJTWQmz2iS/hKVAY7TsIon7469wQd9AswhTdqL+PMQ7
k0/mfwbrbDtYPqSfxuINELR9zDcEPUh8HlUAoPBHEp4bCuUN14xka9h2l721lMzW1SpjGikzPEeM
bGUtg3gJHyVDE/5fk1BBZYLV7Ung32n0NMA2f/xLvXyMpLhprCE+4QnTKCXjKDx8TPOh/Xf1j90Z
B+kyrTNUhYpWo8U3E1V2PCS5cDWsSpt9JRjuH15uj9E6TtjVHMg0SjZlBykYqPeiFFAdgGETDbOD
3DIKmh0Tm9B3wgc/kvSppCljfS1m7IEsNzxwgdWEMotgaGfLYXmOMeHcXVN1IK+pR0C6ndixSV8Q
Oeld6JvSArWR+1oiVHE8r/NhE+OEhRV7/9c7CRwQBfZai0g33lrxAWZUOq/aXVfv9AKZw6zOy7cP
uqYhU7o7P1Ti0S5O7LGEM/ZoFE7buPGCd66u/C7PIW2rw34qTSpvi90VfVCikj+q6YiPUX1p2/CF
kJ4pqM6X2Q9rPQcUa/ZyH+Rc+PuuH1XM0wJm2Fx3Q9b3TU4OSvRVdnycYC76Yt9ngN+imCbQuCaa
zPq+tRvbOP2+ZJRIBEM6YzFQzwRDSPd/1G+JWmEzSWHHers6yukXsi6jlPW8ZtOAYJ5aWgRXmIXi
KScF66SJv4G5rDU/l0tw6k0CfVZqutUbyBzBELqncUoJ+/buCAyzPux72iIsXY+6/9ikLnOHOOou
YwccPWFmgPpyjYbOyjd/JCnOrOqm+ch106N2ScH8wZqOVT3Nb8wNtynooiw1YaNr6HZD8dCas1HO
7bv8dEgQdwxPGN7jwgRfIk5IOblNBYIUWtOo4Zn6mJTvQi4ZeKKzKSKnG1j7TkGJXj+6KqLzUExM
hFbdszI8P9nE9a8+spwitEVuxSTsbHUgCvKoUNtxMsMiOUshE0KMbME/0oidAfV1foGkeyKccoyj
WoYFxhJ8HjJEMkCCzJrC6na0ZfFgPnk3aWWCLWl9CY33id/QQdKSTAMmXqtH4ypBJOT9E47aOrcz
GZ1+99EMz7kFpCeZNMBJwYfswpjhXboBzuCOk1XhiN8RzujSFtMxevjZGLExW3tD2NDPgMLgZ8Pa
QU8xHMqHeWT+AX4BaZ1D5XrqGNV765sdKSk2MmfTziWYAwqNmc6lOCFnHben0+3rVxyTpVF8ztsO
d0GgvZ4Ib1C/EOnzSxj7kfIPLVliv+ozENXxk0MmcdYS4GIF4vJI5pJOCZ3rJssFNCnlR0ogHQdK
l7H5ZFi8uOsgX7OjJqb3zAbnnxn87lOUcXe5ySjbYYiULxMSCR1ByjS4k2LK+KVLf+2pnq0AJIHq
n76j9/Nh0MhEIDwz88Gz+BvQyxIo8sFkjNPIRtPC9MxZEziDgVYzYW7JNmre/9pzmOMOw9WU8/6G
lOrDJl2eOX9mtmP5AhNUdHhvnAksCwVXAaGNKmSb2tldIRdyxFekK3jfIerA53feu+YwyDfzKYYo
6XfRSiVNvSP6XJJBZlB1cRDj9/oiuj0lsP68gDcXKsBPnKPLjgRUgMEzSF87icpHVs6iPVxd1BZx
E8Vx5FCZ+F1sKmz0pBXqXaeNUb7l1u9slRnIveGepStr4MK6zF7WUNPuwqj/esX2Y/hA0ZQtPl2h
G3vnq0taIbNNw9oSpkWeJ5YeXHFpOsuyMyiCg+KWYDgtskhXwuL5hJFFE9G/yNe22wboQ74Etg86
ysFJpSBxmq6ExdaJYqxO80k+a9fPlLqC681bKSYYbDj+8ypXpCUS93xUk++LGAHLHzqiAQGBcRQl
zPSFDlVWakXvuQbcgGMEm0WTX5OeUmfkXiKdp4OypXx5ffS/7Jq1VRXaiIx1uv9v35wiQM5YktR4
ll+ia4rHiGLYZP7j9vNhRuGObABDkSl6M5sYMclpR70moAIsavvW/NKyW7dC+ogvMzZTHuXsn+iN
uk8dAh5AXqizFExCFLuZ8QxbgJNjjmCAv7lhnbY9m2M56bsWnA1r46Te/hjpHFC6rJn0TsvBiao1
hOpae+5LTlhCI5h05EwePYSN6+7zP5iQr7oYmgFgbnhuYwGd8RmJD5hBqBjqLzbbHi6C42lD7tMd
wRx4cxkvK8K5nWFsWU7PLTwr1TqmynemZfVOA52Fni80fwsiKUvxYSBOHd4v7o+RSkKyfEXKM634
MGXYRwJKWn0KKaGuwQJKoUHdPv+0Y+Kw5jYPCuspmMlAyMmrGhOyGHSVP6+gXYf9EikXDXp2PV/R
XeVpXxa2UCh2+DooWGklU8iAAqGsFaVh0ueWusPBZ6bqn7b7SIxSHxZARM/vf4qooRA7c4COTj2c
O4eFdw0K6bpe2l0xHnuCM1HRmcOLGVFRbb+pICMEy8VoTNfgTfP7XblhJgjkYoOryoW5VQkkqKaV
yOiq9ABiH9jlCcQdkAWZFJo6vTY59O7Id8mGmszvQujlP9P5aVcMb7R963QkXZDDc9vO0MM2uMNv
z1/hg7bLPr+xPlbPjQARv3c/T3JD/BlZ1anDdz6MverBJz+GuhJuYMfdiR3ProO2JxFZsOXic+8Z
SR3GW0unWQqjN2mWuaxLvH/WbSfTn8ExRTmNZyRxhcNLKYJYWaqaoaHf1IsStgnPwXFnjMQSeXfz
htoCQ7Lp21x4/Bzjzhfy8TtBgcdPOxkLxyIxNzfr/fmSl1nZN8mCwXBHq5RdwBfmhV8Al3SdGeZM
wnMkbq8QNsZQXRWxvLPtyTC83pLmwYxUQESLBmzOpgJenQ7V+uiznW4uXhIDlVuzmH2tQ7tjIb/j
Sv1p/QDKkPTPX2ESSdMGHfkxTKI6tad+D8rDpJCv+qMaLLeXOTHmj1zucqE4Cny4ujHMUSjC63/K
dwt5sAn14xFLfcs+wlcMmn5530/uyzK18M7vN/ajKZ95bhU7R0guQMBK7TWg5BjZqWOqCS0+NU4g
Vv4pLpBUSAOWswxjE8lCk+8O4LqQpHfVN5ojQRcIWJgY1RN4rSi0+Ly6NZP335G2f/0YaPd8RVPS
oe7NgnwmiSofMjNJdUAiIKFcHCcj2LixcTs+fzgyRbQvabHUf/+5fwWOvxrKuxPsS+8/DVDX0Vsp
fHDdDD1nw2PMuEzRNwvMr9neotdIrk4kJdLuEHcMKdtVjlHHaF74etUrG60YbO+ACG47582cptdw
qgyDtOEESoUBOzElRjSpDTyZFucfQCRC4/OBluokOvD+0oAPLX6zdpGzCxIDHFRQQN1gna+bVlz8
1XK8PdT0HQLbeBSz1DMlGFKsP9o65pMlXrqIwXdXXrDvd5mV2CtlEfSvXLdQGybVfFcfKpcMsRi4
S1gINHEtFwCsSA6graKnXYvZx/XgO00eKL8CsberGjfYZS8NistUaUkcAyKrBnB47/jlAg2bP7ak
FLZ3R/UPmOtBroILfZIzvZUUiL6wHpFTnWiOip8Rk5Nsb1TgrKwdcoMdb8/Pkp5EEmFYbm5Ziz7s
ZUObpwwImuPYW65K23s/pGsFSBgFw+aaP5aUIOb28UDAmc2UoDFhsrMqr5SpBII1lxEv5nXIA+Ow
6dLWE8wpOYZYQQFHVo/NbsQngFIDLfiDmRUHf+t4tqH2rN0SQjysywYl0ToiaeSxiZbfUl+GZdHg
Nxk9dv8Y0cEkSRTT0ocNCetlbKPwaPZYecQkMJYlH+Vw+UJA2nNrKTttNOlGrN8tqiYB/5UwIpH0
LjknzBuyKc5oVOnDYDZAAySAcW3xjzBalsQZUzuTAPFSvrIFxyK/N0R1KbZi04Fxkw+UgIPjxdUv
camyR+w3T+ryP/4XJkOEmLvj5vjtHT3N6+tQHiHnxp8nNsM+up1V3KHjknAk+6XkzDpc3K+aHKy3
tB0SVfRYbg07Lv5DrPWdHpAxCEOzPPhAS82SYlsr+CLCKoySXLHtVQUuQXLSda+YX8j2zNLcVi6y
cMDwb/UeW6O0w1aD32h/I4T3KBaFcaNea7uTY/k74B/V9z5GMVotvpViZgbQWthhbf4n3748t5gB
n/89NVok+D3GMaYpsMwwn9WG4GXrAtH/yr+p817SE96a6CkkF5JS6nNEW/EJckmfIfa0UogBc/UU
hH0IaqRZ6k0S5DjdlH26gIsf6/HRys65zxT3q6pKuWR+eRoGbPysgnSEZNE96Tfbr2cW0/76dagV
T8Q3Bkv+BSZzeMkpKRssifASxdCJg7ihrFZ6o9awOAm30ubgZkVAs86cGJbMsJAI74cZt5zoyyyx
auNyZ/Tnns7eRZPKX7SJhGnL5z+5BvvHOMlEGudetW2YCUL0rFMTc+O4uNEm2yWv7AGXPaZUp5hJ
HWaFkmPDAkEHvIE3ctQGmoGyLN1cxDutHrH3tgE2+KcQKWgzEGrhw4XbISyp/O0vw4p0+SeooRVP
h35xUClucn6qzWiX9Xg0tvcPNg5A5lmD57HdQgG4ZBESt1z2ER86Upg/9mn15kOzb1tzK7asBqrn
1VtAAuzA5r5eSqzY/6Cfl4aFTOGesvwA1t+4vSHFtit4sDtuj8b32NGDUgGggIKkm2OmCV7CvQMf
rFXkqLjsoYrD7F0IqcNCEKhToSoO5EnV6WDFtrlla9rJUEvH/B1McoDcSpBg8Vif5/lJqwOqfKLC
XGX/SBlw2Dbox3LyaE4/H32D9UQPDRzkR2NCpWnmYUR1phoqmVP8Bu4B7+IDyKWA8xfDm4YQbkIr
FSAfk707pGAUQmakarM7qg6Y8bj9yCiZ+JDFTb+5rEr8TTTdajdhmJ5FpUpeqK57DpxffAbkOyA6
uUhSgXgd08RF03FU1PYw2GEj+2mjDckSidaPtI0Z8OfJ2GmzuUx3tXyxv9giEqDXBjAcenVxpGf2
7SZJGdCH+0VKE21vVSqSm0y2v17KOJwmBHvHEhdX25/qdHZeqYkpQO41UVuW+SokoKcAGlrN2yN0
ixoja5AKdQ7OtvNRTgCVTHeA14QBDRSOmDXmC/ghfe8zOhxFzIsMy1DHG03II4TIO7zz03X/oPLI
kx1coqBShr0AlsIvg+O6rOciyM9Gx3ZkHTJN9tsp+eYt/2KRLJc7vvm1vVIal1OfzgSOZwByneB5
Sx3Vmw464ovUktivNXemQ/4OMhADZUDq48Akgu1YrKfgSVs5bwEFjyiPUES+Tcm+4fFiKPbalmsK
noDb0IvMwN878nD9xlNDHGjkkK9NK+EK/ebGxECOOju/ukwpCVAwpvEgyDcCsaF3DVjo4qeh/WRa
KHYMCIPDygaoupacX4b+DgfJnj55eTEMIFGE+g/y9TtZ9EbSyWjjiHpLyuRhfBfKaEjAXR0GN0zT
SJMqniBtMxMNZVpdU8XNOWmta8gdBN0q3AlLs0r1Gk48OZjerjH1XI9h39zXoKnyi4PiUf9kgUmx
Yw53YAIHOWCGvHvMALgfAfm+xkWQ7KeUsWTHSH/DX5z+CA/+VGL31YeS2jWnHT0jPQcd5/mObK+n
la34lqrcVs41DNuo/MzihNRF9ESmftysWW9lwzoPOlpuam7TTwMsTXIsEDJRCZN17VEpQjB3hUpg
98yM8eYW96Hz6oZMdatBLz9WsrJzM+wIl46qR2g5gx9DDHV8rngf1mpr8sDJIFHcz6MYCv6HwKKY
HHVVd2aTlpuFGv0TIw4WRXIJBUcw0uqzYg9DYC3WKtO+K9BLIu8eaPRhX+M61A6XQgr3k9z3JwMf
z9MXQZJ81xH8QMHwQLlj9i5TIIuD1jKmKHsowP6r/g9JLkgaRetZumWTtCilFdgQRhqBXWygmuly
TyeArpClclT/Y16YcGJDR1H5c6yKSQinbOnYe1UftUAtm0WfEB+lBySRGGZTLEx8r5RDb0iYq+Nx
bepCtkv2CPk4TJqW9HwxCRNX/2v+0O4un4Dm0A5IWOx1VXbF+AwtO4rSK7JnKmMTRXsnKyN+J9U7
Ey3Amy0b2p+L6JY2pRlS4rNOvnKgmNTRCMVeNDF65cqOQi67ZVTuolFVU1SGdmjfvuwdWORO5Cs9
JzksCm8RJQioRX0voV67JIWQEoAzzzIkKtPFM2zkwZf/Nr9n0gx/K68pTv9DUzcnpcRfPpVIRX4a
UebdjpKVWduTY+5RhSOlzfv+6P9c8BZmO1feCVHrysuJ7WSTFe5mNXydzZfGZk731klPXklPyU45
8D4kA71WWG2dXaLYfcpZbkUFDmjppL9Vtj8fPQyqeFqqCLL8pZqMlB/S9J9dTSJvRU4x6OakJzls
+ynXf8auffDCNseWb+yZ/CLIAhF3zWvF/2eK4nP4T1qjfVoCJycZnqrIyf3ZeipBThKtj5NWHxcd
L3uxvHZ7v8qL1aeNZmP8FCqfg18B5dwQEAoQcJykjlhKpAlomvSu/tT4TYx4YcCMKUIoJ3jxNAA4
S8C7jm/WOES02JctEyFZeSVISVQ/zXzQ7QTttTxCw65m5dBF994CpbjtuUtQCuNd+Z9DsjeCvDmg
M+G4RnkPhN/kNk2FF56lCUHgtyeH6oVYnWOtuedqRqFVKerr69te/YC0JBf69crgvrRUmWyoVgHv
CwJPG4pL2QfKBOOIVDZEPnq7ZIKJLFp8bWCLMTmx8u0LnoJgP96qrTvpJT4AukhvMAMKn4kZkp2/
UtNiEHD9VxcF61eGVkKkGRXFtoFye4MB68l1TYPffv0XE6PyScFjroT05kc4Zwh/UFHNXVIjSU7U
mQMGEIRjlqNd8oB3LLvGD+XmJ2rl5Fir04TgGLQudu33syp5x6RR4xEsiBFcluNLKvJGz0Rznklk
Rrxsu+Dyhuon3cNQAN3S9CQy2PQCvtxUJxT5WzHK/u5xa1lf9aBY7a1KRvUcgV1+5V8Q/tgb9PSz
H0KKdtTPaGE4L8R2z9bTKlM/5oWc4ZDAbyCRyQoxfJ0gmPJIfqhfO9Sz9ASO6++pXegRdAGifvOt
+00cGAS5OlS9WcSTQosdOytXoBuVCJzKEH1lDgLnKb+ixFWwz3eClKxjpun6LFljtYYuHSKer2rF
TKYWq1SKetY/4FVGDrILLz1bbclBYcjkdw9yFW7IIRao7/UBj3vqxkxE8S4PW+orcQ4Yqt7Zcpzr
xwU1bnYFQNi04Uk4HcjwGHXX+G9GdYBKELTpHiWEUyTB/Ejo/rt5r0J9iIqaSclY326i658lxkxF
UfVGB9fWXUE6W63DUpBd/CcZ4wMq6MaVEBQ5qMxTi7IgcWdbYksbHuu21lBFbkClWZ1oMDPWcDDW
mue9V5LdyAsIKa7yktZo/S8R71ku6Mkgp5PV8kboQHABrrqlduwhGiAHgmV/qF0MTqjPjDYMVuxt
0AzeaFQqOTCc37ChWrwp0pGDhHWDQJUWMr4QgnkLjUZGQ/sqLFPNZbFYBnYkLb5afK4vEKBVbZON
UZBGChRHPrEHYXhsmfucG+39oHzAOyEpd9VUlqxZJMmEKs4CCLY2Cm3b9l7Njy9Sj7r958I3FdnW
3KluIKfoRAmC0VLit0T1OeXYmsiPtpE1jhGucS+MeEbRf6NiZUgoXeEe54AoRp5zOIjN9IjPrehb
ymigh5vp6VR5cKFdOULmOhGNAFC8aDdUdMsQ6fiXTMtIJIwd+n522eBlbJj3Zb2tn8xK0W9qTre3
xiyYQN+0YsJa4LGFlnd6tkq1ZUHvTyR9fTixY+g2zpXe/47atPtESVrt92VRTbqfmItrFBbMrGUM
RzMrcTiy4LopjGwecQGZDZEdEQKbQ6NmGO+zyqO85kZo8R3g/U4JvjhRtHj7Bpzmczwp2I0M8C2/
610NlzwTrYRzGELcsjwRH4PoZrf7xU/ZA4yKATy6ZF7mCzKpIz1K+Fs5PRLHxbXBPESDRB/6gfM2
fZz0HPXqmklY4Pb3774gQKTvo3AP7XDOcy9ESFbmWynWRT+392HuJyIv+UKt6OtMiCQHW/G4gkqL
451sfLg5/3oLJ3/r/DDx08tvvLOw7cEoL67Ky4ZmWd1+5b9pqQe3oXH5/s/yzjyx7oAE7Q7I4Hw1
fpMTVFH1C5EL0fYNJaKhUbaNufu/2vY7YvD9p8tj7HpsLfUHNkE/fCvg1mzjMGxtpvGWuzPww87F
bkSZEDqCHaw9QKoPEeTSX4Aq8Kq3pkM4E5aGATrchSgk4+U9s4PE1pMBWxBAA4yZmhdGNcH0Dsjy
np66VnDtRx+cFv1RvpJWwas9bc8SB7uvIU7WmlZZZOG58EWxzmHOTv7UZ3VdhPwvK6pm3XAtx9tt
WvdQxeTPYOTlBF8tb3hl/gOqj1y9hv+bd3efH9AcED3xdbDb14d1zGq5DdjwaNPOFmE+0WTGhHMC
wC836sf58MIEwx3B30rS86SH9OQ2K+jpA7e5AmUxoDB8l4D1wz7AcEsbfvZFtM/QI4ruHN2BG6Id
beZjc5zrR3vi7vZMVilPaLbIf+lVJIcv0lQ1yvmMwSIQE75R91FguuQPnvwdF+CzYo9w30Rgd6rc
k+oWoinkednDNVuUSEYnmOcVOshJFuXBRZQIYTaL2dzlJkjSrMU1D5R2zbBLE1JWxZ5o9Orn7P5a
u2rSG4OtxVVh1f+V7BH1ZnY4EpCn9eb2dxDHeB5iXDFbDdqN3MENF0uQ5+ZtxmCvgzBKUbVq2KuM
sdJ1bqB5NSy+9uv2vKAEdwPXO9sbiA+g0ncBllnF0Vt6DjWTl9BYr5M4HJl0D6YJjrnCmBfkZMpY
CjBObER7poFTqXn+iMBwLIX94brZx7md/sWed3EiB0swM2weaMrEIF1vpXbauAr1E9GcJCr2JMMh
bO3U0YF902gIXYtrSTzdKXcxsAUKDML1bhSniFY6H+m2dZ5snmrhJfsuW3/dLqsZY1a0pd/u8HMr
8yUC0vXy14ByhB5VdAiSj/vwZmRQtBTigqGwlbyoIxEIT44RaoCWq6E3UrdYYbw0Y2MUltgJueBE
AtGXW1orcWXUQCsXC5LIEAQ3JI51g0nx/DJ7xiDfL69hZdLyFEqny8buGHiWF+Wqk3edTSEi1EH8
FY8ioOWWBHCF5KykGEFXBR8OEWw4eILHc2fQvTycHyTcIvjcUfz0ULvx62mN8KJAbadREmaAEwHA
m6J320SDlF+JJ9sfWtFcmrPtpCLKjg/hIg6LwXRHkOW4tjqYeBku4rMsbBoz3w34NN5wFXkRfWtb
het4dLBWnjcQQQ0lyqoXQayWAUsJdwtgTd73cvfzEdmCWMZsDetZW+Ptwha30eaElk1gCRnj9CVz
+YFs+Ichdhyf8He3s5tueITXxIoj+SG0YpLjUN/F5KGB+I8RDL0t2qP2NA/wDJkeB1iKz4PbVvx+
A/5ivcQGIJDpVMiTcti+OuLsPfXLaMVpDkKI1cHUs+MBJywolX/56dDa3G6Ci7DJV+fG17HfoiFE
51ubJRIJ2kMIgVWGmxMGet+XKtNf403Iv1gaSwZBv91UFaAyQ9S8AvesGQ1HHTFlzQW+8xb/BI0G
A2KxiHFVcC2tZzRUN+aN+YwiFcsTPI8hWK4aOC4kkYT3YpeJXMWW4VwE902g5+epi72XNgoZlzxz
hLBnVg7zEgQ+aryrxV9AZH+L2YhHZxe/5wTkyblHzCFUz3+z4aVgw6DoaE9hFCu9b4eLSblzqlSG
SO2RDL/isAt8sM2vkUuuSHMGYh87fjkoyz9SEAyVWeHrm7qfYfRHiMIcKPxhpB3PVrehX2LuO+zt
iVpXY/rtd7a/k9UOCuR9a/sPY94StCkl5voZb2C8el/ChLyvYjWeV/sNMS4drCaUj8LrQJ01/cUl
EGZS4qCvz9UiQyxzLIv361LgXJRBjMCtoMId6egt/Ofhif2/MRL1d7CvtA4Foxqd/jyayPXKbtQs
c8GiLNt332k0gCHd0vkw0c+ugHtJleJBnX8VwE3C3+gkzvcNf7BOZ3W2oMmLwIatKBRnSLtKLTvO
YmVN9jij0Qupt9tcPi5CNFaW08fbrlry00Q4dwle9QpUAGaUAJJXe2mekw9AApo831UnTwlaBGo6
KiMAyxdr4XrSPPhIUJAFLo8kseo4IO1ETRC7u+sobU1ZhZUCr+Q1EwTouTj4d5bQ6f2+zsRgb17c
/f8T5oMfmMbqVhFDHvLZ5xbQ91UDDpANzdQPzxyX3ODmhdJdAizhfL/mr3sjv0wgWpPKxX3UOaMJ
495HluPIpaPNjVyla/yJrx7ybY1V4w6fWhprtV3vZmzZcBioAACf+Ay/PrsAFwiQwrpqKdVjaLTU
ZA9An1daP5/LOCCkl4g9ezikf19PFMVoegf/6RQQjvq3+qls7UgZiNjVogtKXldxMkMsdXnoRTZQ
pRVAUdlEo53RsMEsvZjuw5pf1LIJW/zP8QwOi6Em63itHxMKjRRJA9pBdoahMVcG9l5cXoL2PCaW
/3xe3PbfXOx0RZfoe4D4yTBA3eAqJ8ZGdyqfwrz7CU+DjtLf4kv9cHtvOHawqNSPO42SvVbeq77u
beVwAUoHD1imrWlRxka13t5Hs+Eua+4tI4XEXoU/08IEQJkAzsjeLGTqM4egQMNrVP4PqxjRqO83
0iu7CWqdDNPkemguBirckvv7PMY1WxJSIOlxOREE3J2YHT9+ohB5wi4XxjHx0xsyah9+C4je/Dcx
z7w+4oWNIIJT4l1lD2bu3tOY5jikaU5BqHZ3IckWdprxysVGQlWlBtTSrwaFnXcgu9wFSNyYel5v
QgAJiPghocGcuUggJi9Y1WUX+enN2O3O6hHNzNFhHzbJ4us38Mc1HsRAvSkjx5SM42lr6B4WPqAc
kexGiDwkLG3NPx+t6+dMmzYOEwbf0shHYlmSDAuiUm/6pudPQWK4oDNzeL09+XmYJYuCJhYUwnNy
ebeFlYpzpsfqHbHucsCgvphLB3QyVRxPPfH1hm+OlWcRCVPDNgj8D5L+L6BePBTO9Z+NsHCl+n5J
YWBxw5OPqd+6kB2tt7rQgAEO2NDEw4xS/OH359N4TMRYw6HSutmWtzl+Uk4hLZ+k4ZL7ZeYsliL0
O7WWHqkhXpyDW/f/LSJufO2DEXb3Ag8gxrkTixtQAN2SBnO9OX6O+KJGK0+PFngMCy2LFDBeAvG0
h8ebwWAu3vYTyORlNIlVuuH+bKbWYK5I5rn7dYiuLUCawxU5kS4YAbtPXgzQHn/m6KRMQLgtLmWA
gbmFV7dINr+U0oSh58eNteHW4X/ETbGtvt2QI+AaGeoxBXRhtyBhg5j+jGgPDXzqu2eoJi/UQTzv
dFb3NEgxNA4Eo9ubY75FexU4aOLbWi0J11Z96uOLJZ9JV8DTMHXq3oBzLls+Co4PgVfrq7mnvxhB
rZT7KOeNRTgZPP9/gOqzBOAxgDC2e/wKTapiKykZNbHmlCsekAHgk3nhYhnwwXrLhRgz9rJ/cF/H
lSeoIy2jv/fylKDvMWVQDCPlEju0SzrnEAOoAEXSAeSBRgUkUxubBexMYq7/pg9U4b48k4JYTAev
+Qk7o6wTQfvVmIy4fA0qw8E/LAw3vb/MXbG0uVH2RgDh5cGgNZWLGplzDHz9GLLDGNBi7JncTgqG
77jGZd7TRyZMwmG+9NX0Hk87fJw0oJ4YUsKWpgRTpo/wOjOYZKuxNUNUCM3HKguDQmN1lZYIkSCS
rMWMZioYYO43eQP93GpX6dGD/SID31I73ucbEu6GDyfGm4hU9bN42agInOETj0pA24Sasc7PZIhI
t6yNR92NDZadpwnMbjIeoHgy/lrr63bWAfWUPQ7lPqw5SLPugQNo3Fc7E49ev9urkYemErGMudfr
I1bZyb75KQoIWie7Rmj7CyUgFvWY90qogMYLDU9oKcSWghM1vpVQkpLd/B5oE9XFV4jgclfBYfSi
2HbyA/DoqjZ5frjRauOrbtKrNxn9eQNqF6qjz32xseJzPh10NU6hvB8RnkDryDBYC84oyqh6OXOp
syM74PXxYjTt++QIuTcw8pHwV2o/pPlGzWIpawYrkaFtf7/0Zk4yFpQ6AWhFZXLXCg3RrA1i+yCr
bWBVCJemHzpbo1mfUm6Bjcg9MPCHySs8cImJh+dhbfFqBfdGcsydfXNnhCrsdKXoFM3l8d+7+WOD
PiLcIOljDcPaPj7PKuWE5kJvY0qs+KtkR1F3Sglqw4+TD1cscW4ewKiFWMyRFQQPxtCEliBAAo25
To2LUuqK8/1MR20eYL/8pQwDVerFikHlB26/X30PxbUD0n0pJsxWv8eKTDBHZCxK3Ojm9CEsmKuL
rcknk8Nb2zul7udy4KATH6s1SXDs7Kyu3P0hUkMSbft4LhxF2p+GnqjGhxp/8UNgEWw47GQ86V5g
veOhmoiK78WaeYfi1AogOQxbI5kJKQAhS6f0zI9GIIn8f2Y1D7oys8QeZjC6vOtH3ev20kpnEETL
rM8Ae68rXwEOGCfGSNrdU0XiER+UiVekgy9GJuJVTLms03xG0f2eJaAiOsyFHVi/TBA0EZNQJroa
If49EpGdZy7aggR7udS+bC6Dewr0eBgtIlupwb1ngN5+AKCzrghGW3AlJdLpe7spHaFD7cS0jCVW
/fuMy/xWpUp44ZnAY4PhTCJIh/jzWJMTVEndSIZ6VezH0jaiGwzHknSFQTFOMQK8SAryar9wgrIk
GY2Paj5cN9GqqhAVVtdP0i2/CR/e/UQfj2Ty2iHmQdfBi8V9p5lCjNIsnDuIJCTc3DKcmXoLxvqb
uH6wyGdSpKyIAYXzW+sRgU7XsBo6Y+HS6Lpuyw9b44gpsunt9oQTDCJW+uheGgfWGV3eooZaUkKq
AHHmINFQs1kdmOJTBmrJ4t3Bfmh6/dIeySA5A8ubw7EX+hLe7+sHuj9fkDr3J9N+f8TS/1qwqiZM
UE1Y47LkIstfCGYBayxU5carlvcM3jm6VHnf0A/7AS0qP1jF1mh9hrtHu8Su0j/MGgkDTB7so1aK
tprjAA5kji6lLsb6sZpV+9+NrvxRRwshYjrvxJO6F+O81++anSQrsouaHvHDm6N9qHSOwOWOnW5w
q5mhAz0BGU/rW9O8nolmcyPGKA09vFVUbC6uNYz7FzeFQVpjPIzf4C7WaV6HQJXj7cd1gcBPJCYa
HFHYmJR3LdQ6yKVfQvxo6C73ZrTpsjiVwV0WA3nISZ2tf0yYwPQCbm8AR3K8aYDWYFD5E8LOKAQK
6Yqzm1EtmTmfmwdn67Wbx2HKCWVQzzg0xAa/PdKq1xAzuZJh3CqGiqgSffgfx/d9XCq7mpvHit0d
lzyozfs9PYGqhkep+apmaXubqs9ra/tKwetW/ZTj3VSdtNOR1nz4E00OUcO5JTDIjFUv3kiP3ueQ
LtwMAyMpCQ9Vwcu+/tNAMWdWa4ezocgz+Zsc6OoV1bjoFc6joA06m+2BHGBZNXa8rsvJw1A3qz8Z
6Wrjwgk9jnai6dlqKNtYSO5260/4gQuzpabc2wmXSY7G50dURJRxCCIPM/NcinZh3kV8tv6g4+NW
GrPW63qDtdAojb3p3bNGH7J3nSUS30WuYm6699t6Rp6tPs60c32zgmiV07oieg5Gd2l/jS/q0Bs6
8ZMXa0jDsMb61YAHj0FkbmYcm/NoTMao6Tky/kxGWInO1qzaF1sqS6bQrKD7bJjAUK3+9xakFTqW
ElqlsOGnN1zJx5G9zciRdlXfF4enots6B1FJhT03urULZY7Q6+Lxu08YlzJCBd37q+rw3WDjuVkN
3UFCHL3vF9TL1llE0PIGqI8gdTfWdhgde61RpNDWQXQOtf3d2jn7uk/ZgOgqcBQklp1auauBBj3M
EMeQVvynLavgL/PK5iMj9Qn8s3lhWWYxepdndcx5tIIyG+GDtk/HDZFVI5klKLm7al3OdI4WJ0M9
KlYoDMsatu3MPNY6yVOMwIyF2UmgKEjNDHiqK587cEvowMvxu7QW/Vv3/38DvHQGBEZw6DJMwqtY
Ldo/qytQlbPEVp0XyUF4aWeVJEH7vQOIP72f0ybdp4glli5h6IV7VmBJ84ogFu+/EpVdFD6QXYBe
ia4/PpOW8ojpRqMTAcnqifSLume+C8MOGkDSk8hfWpgEbgO7jA0QqRMxtyAIIObxwlCDJVDbWjzX
G5y7CGhvZ6UwstZUj5EK98Eq2mY3TbwPQOQtJW/MG0UIC7GN9efgb5QWc9nqOpsF5WO8oNZQDwMP
Q59y+fkyALd7kv0Dyue62PUxxKqnn8F++Trnco4dpGggrXt0GpEWZNqv/ZG6oyOnYXG/C1Vs8OtP
S3g/ENVT0rj+a0er193cWBrYHePJTimEflspvOmPk4rgtMlgo0mFi4S7SwirsOxti2OmrrFQNyP0
IyI4xM8R4QTEUQJ12wquYrOqJ9YXvAfuvUgeQMM3OlHTE/VubuSiL69f7l3dM4CeKd84twq7mMgh
5/T6bsVzYQ2llV9fNG1fMPuEWRVyY+RwoElCHStZIRj8fDN0OaELOSjqahasQOK3+9K33qMOww9F
HS5QO1JdlpJ0YTcKdJIGloeKo0foF9ay6vRW/ofl4QrzbVOlCA8htb4uaj/EUsg+hoA55y2xYAUT
1Fz7ZiUUFc+q49J9MqnuxCa1mBo/Iv4in536LUf3PrnaKsqiwqEEBwirt26QBCivjJ1TGVMxPnv7
po6JN5Z5h/Xhx1dOE4VsTSllm1MYD4z5D4oPUltkMUTS55sGLIMRSTaME2NalYl37G9KQjzVPCdG
WlY/wER5ZCtCcmZKWRhIDVR0HDwRIZnWnI+vrmCanHFbWIVWLX50xwkqEsswovryqAq2DKKq1IAR
uIjm+pFy0XfB1pceMX+wRTcMjpGpIQYlTlefumdgPcZa+w9MfkQ9immhXBNMkuN98ky+wjwdNExu
WLJS14Tu1inwSVRvwmReFJC/uy4tC83tHN5QYsH1YMAtxP8gaWif+NmrqqA7bQ8W8ZcaECvcSrTz
Eb1FQ6DM17DbuGiFWN8oogc8ZKps6zidFb2ZGBJW0IcVEN6RrNSAHBLCKo9omkqeVpwG5eL1TFtK
No+P4Tf61+scyMnErUEeG96ra2CqvLcjxwiqS7ksxBYOAujrtknYr66RfV+ocwG5YSggWHrXvACX
eBVQbA0dULvtJOD3wiqVKdo3vF5iDliHsvYNAlzohm0oOBYDKajymFRE4yX5eeR4uZ5MfEOFVEkM
YvGeAIz+Daa4m7BKwLVy4HLwYEeZ7JuHXKoCnS5rKsCjAc2vCfLGIawx8ZWP13qEAuf0eemyNxuT
w7SUXavK3YCfI31pv3Sl6DJpGyRKoyM5gShUVwwsgJ6O9cyrIFCraO+be2IVR6yvRnY+JW9jSr8j
dtC9LhQ027UjBA8EBk7+PFP/iwTY0IDTZePIWblQUuIMrPB24c30MAwWsXURWaMyuNCm3L18XVDF
NZK8qtQ0ulbnrsKQUX49MtrMWGOnhOguSXnBe2YdlMIwg/wjP9zZyjwooAz7dsUOw1m/numG0AxP
IMnQAuylNFvsGbhXIuXZJt/gimWPUlLgiYtqWBCOATowSVAzFVRyOT5up1caR8ysu+yzXXzjMnHr
dUm5+AeDh72p9BZm7huBCcXvVPF9Ua5OKkjqNCIWKBAkBAonGSCQtfzrykrX7iAX5paVQ8QJea0J
aIGbfVm+uqqzc91AWbNr75PjtyTXGGloLkTjwLvVSNuiz8DrjySpty5I6V6jglQL6l+Iqn81gG3q
LChvF82cN4gwrkhsHpi1chJt+PW/2CdahxRMYpeQpRiiKyyNh9RqFqGnI4p6++/kcJwWFsbooYC9
FxSB2vSGixAlTkIEEOIaKfYKRi5EBNAFvag61gGkXJapP1nDpdbUFlKIRCeoj8friWnPAYVR2Lud
aNrQj3m/y9pOthnZNje/+QPgsP0zkxyG0gExgTM0gMX6YWxV9HOx3mlHKTylOk/po1T3Xu9eN/n0
/7+FRNcBsPMxIJ1/VUpw5Er4MZRpwAmriRvTSJQ8RIt/6X7ySKSecx7RmqzLh+2lTTHNoW7bPCL4
sQmQ1V4Npf6TZ6cXBNvtPAdeHXvJswUWeatqinrnDb/4+EZ/+IjvHhfYHQRNzeCqKjAay9bIWkza
wW9o2Y5HbbDuAbM+RbGwWRzcbUyazSIlXrySMUWVQAcgncpBeUQgccYLjhq1rroC3BLfv//UY8yq
i3Me3YsQJ0LZZQXIAD3BfGLKW2rYC16cEj9/Z2NWYKJTTE/IbVo+oCC8pxuiEeIn5zXxlN8roQ7Q
m8V11cDisUOD8fnOMNSbj0i4azLXiRKEkYUlVzFOvJjkn3b+cPpd569lfj23F4eAHvKsSoyN3TI4
qadAGn1DvnacMEZG/CC4sxEZeTu3BbLUEISWVu9FkqNPfuqfL0JVQ2gCTExP5CavdQQsFqQy01yX
1GAWWXGdSkygM4HEr2JtTd15CGMTKOf/ZzqL55ZRH9eJEwvgB13vMAQemLL/OTZKZkW+09NiNO0I
Rstm1OncS2N1xvot+Tzq5VSWsxWyXe9vqvxzKZwj9ApqbavVdkarVTInMTqr+XepEdn4v8jWpD+w
8/H/wE3Fo3jYC8CzEZ35u1KOC2eq6DVnPTXIsDq8fHqiEhuNqrd+5CGw04rCH79W/oC/rJXB6hTr
lXyh+0g17QKtBe71W7Rvg/0lJpoof6IWRxraMnBBti4AvBM0TmAoGrcRzLYIWvALp2QSGIS/Kybo
C4kfYkUG2F/pkfW1cj2d+SPNXKRNL5sznPcBFGO/GFhDi1Za2cbIt0uJR9xzOkJU4/4MP8LAbCPy
X5TR+jBXBZhdcLRVUTEMTXmGC/fbpMVL3BEkA6TrD9pY6KkWJPo98h+rz3GVNuCz+8otosc18geG
pe+3pTGgpdTyacIWDPdZaJQMihyJNEK1WUc4Xuxn5ATeeCFbtZqBbqHhDSscO2di/B6CXb05U111
OAPwJjRe5PHv6tbqx4ilez1Z+n/NRo5ZL6aB/XCr7lRzgA0q+kn4VqAFhehtR39PSsvHCo03DOq3
CavwSgNlXtq1nRWIhrnFZkewIZywI9N3DM6amNRsPF351OpTQLKa2wqbRNH9+8A83NRQHIXu6kcc
ItF77SZdkZWNYQstT9GDKi55PQPzLqmT4NxL8+8duqY9VLOoro2fGzy+k1JdlDdDsAIcNpang/2S
TKl0IJ/bgum/iT4PfKARgB0Wj0OoRsIW6yU7Imch9oL8yjVD0gL/DW7ONSmaEFipT+Jy3pkOQbbO
fVsw0X17NiTvPxlm7SX9X9seDAN10bFjAd+3ah6AwgenWW2MWfuZmuolNgB64k0ZR/0015tCQa5r
RDThtsdQg8H+/yjakQ2bExuDIkSssTBHJgeEfGV96dRPsUORtcoDpA7PRhgyWzfnOmTrEEQlh3cG
P7ClLBs0jbrLKt/ql4jjlifsOnwRUhezGwTBj/df75eGSM2BdsmMM0gfE/vUjMmk2jb8XpuPWUwX
OhVoPRG3r1SzyR7wWTT2wjOqBL+ZKfK6CEWxS4yM9JLhE2WTewqDDZZmeMuizDwzBovm3xwgTqLR
o2wu+frt01EPc0SfsadHb55uB7IGGySv0TSa7SF1XROtJZGB5adfahIoR40Y61q/PXuqBM8Ly7T3
miTX+x9xr3dke2jNTL27sERGmHafFQGHz02VWHGpn+QRMUaUvOX1/KNsgzu2Eq3v5+N6jrxct/nb
hGc0UDy61GPCS5Tjw/Wwc3K2hM0I6f+O24r8gTWcTxfKXtNhbnEJgEFgCLMwBYH8cWrXSVtFlZYF
3bl/F/p8BgHs2WmtNUmoMS3Dikt+awkTmsXcgDdNmy8WBQG7kSJJgYVFVNGxtMou+2ac6bR9PBOX
TcOs1M6suxlEA51oVdDCYPlER2f8jqXJ/J0FpzGxgRt4swXfBqziPuN2AnnYQ/+6Nh6YzXYfzSuo
4dqumT7G7UKDiUsKKuQaw/WONKlBuGtV424FlQHbwSYI2KRag949ZMZY2/keZF/NupeBoP8AU1Ah
tGmamSm7R+DhFxUarIm3pCREi8cz6ZsO0OD+vkPnMT3Ui6bIegnTr8LTOU55EMQT02xSxgF4da0+
8iEibaswjqgG/vkINXEHdhiyukVigH3UOlN0sWYIDkWIEZyM0PEnNUHYJwyfuLwOrG0esH+sTJFF
duw94n6ZaEEjjIoTICk2Y8Tr1wlzsj2r1hXiYFXhsPGVA9x1HFlmGweyC+dqO8IeJ0mmk6vqmOce
mH0+JgiPWIpvybMseTsxq8uAH+GrIKByM3sS5vBu5zlXutaG1ctxYbC6sFIamQ/bUjcZu4FVyuJ9
rr8KL/1GTbzSeOzHFpt2h0fuzcaUe4ymFoqRW0w2vKej6DF+dRpruSjOY2QUGekQypyIJL6ng4aY
gc3UUx0mi2TWQwb3t4RTNjyxeFpGQkvc6szjY6uwJkYytkwJEKfOLuXT5xZiCqtYlIS/lL9y6FUi
ixq4ILgMmxNqAQTmb+kJP2Rs8Bi/3gZ3EzCx+wLbDSAO87ZuiFgYq0/2SamEkhtR9SAx9j+5+L8B
e16Fe6fplnEokLXwxhsm/QxZ8vva+xGZWzJQNpUYn9NSodphWB/aD99F7mRFnmyLcKa22ANfsvnM
YMQwzQxZqVJsaHliZZq0NvYiXMLEVpyT0gADD4d76DkiOzIjdgdfeYub+et0tsuMiIfp9M7yrWek
Y8/5kBRTJZ3E9refVvxxsz93v9u6THkOcdrClkShEGQB/YKCyKIg03moUotEm5szys4gMGotvXTB
jBbY5YwB7xFvCgyw2uaBroF6IIGxQgnhCMcWxF4JHr1DOWud8E8Gha9Qt8jOtAYCoDr9Hs8Zm0DJ
HLP3XR5U/ehjKGaKsla53aeGqsh8fpgeRt0B4ULpBjByLMTmq6k+q5vLzYesasPGZmQX4+oP1Z2w
VVYvIyDvAdFsnG6QgNU32hfdBmBdCHMGzNP6Jm/R2sxTFp6KjAlIidGE7ljcsBqztNfqnMYXI6Pi
PgAK0teJ2kXAm5EGF6nb97DtWuOESv7vdaDfy7UPap/0u5MZo/IX/nEjRvAbvFoPU9kYwcy/DUTC
KXq7LOI7OrA5EJJ/sGLA1EsOw0mL/rZ+M0MFope9v2aiJSI3RXYWknbJkO8TufapdLYf5vzruKSX
uc1O1jeNi5AfBG076hXqzqGH3T0hCSTNPYyhrje9Nb9oPr0E8dmUtYQa0l2Ne/ug9JFRrizn/vY3
O4cthtc6EdmGP8yi5PqqopM3Yv0yRShz96RO2o3Dg1h+tA6TC973cjjH5uA5G962ECEpSvh6nl2E
9tsJK8+QoRoOtElL5Wwh4CXxzbGiSn1M49W7ERciPb8YZEcpne3y7JhpCnERDI7RTQJOYlAZhW0a
EIzrB86/X0JsUK+wrTTcg6UqFPIp7pqnjhXvfFbHP16cQWRUyVRvT5mkiHP5kljLvlWVacI/sM9j
tFcnzz2yo2Ehg1eTp8auT0aD3hOGVjmNDXJP1jaJeB3/X5lNYTTA/Yadtc1IDrLdeR7BOAzSBIzZ
6kfasAlHnO2haRSLH+yGvIV52FxHHAeCLOmIR+9cu3R7w8CvPlwE47FdnWrA0+tqeRmTnFRmA3bk
x8LAZf38SsKt8Y7k7k7oYcxu8NBv75PpRibahHEfo8x/IZ74JvYRGfvIvwcCtnp9vnEoUQc9X+fC
sNoBCtYmXL3DptOn9ghhJOHOOb2bt8d/HoyWqcwnP9/d5TTksJVIkVBPQawsJljQ3Zxmz2lwE/4/
xbmdaKjslADiKU2/N5Nj7Hcy4eebFxZL6F5EEzl3tQ+pR4Vcw7CvnCY689qJsv6piKQNuGtxdX1e
+JOU1CMPQIZyX3/dVDr4ma8pvy4eLY1X4yo/BeDyWW0gfT5eN18bsu5ewGTkfXN/uD9TKd5IO1aS
MBSNsvcPKd7Ypq1DNS88KdotWcSeKt5VyxphpXSKlMdlCzkREdkezYYScW22IgtPG7qKefCwjWcE
wZfURORd+vAD+cqY63igPMg6PSOMMCURQT8/mpmmEOuMlYClAC+B6dXVzyGBandzCjnoas2VImik
M6wZt3Vw9OqObS+Pscq5fGRXHfmjuZ2ZDoBkFTrLppmHQ6WRc5lnpC12UmquqegrmtOx5vtWiQxA
u4L7an70LzBQzzVxluTHXiS4XAUHD20uILEHs/C6uQAPU//dAkCWaw5TapuaOXYVSFqzaUoWeVg7
RzfyINQPQb/xZAkapDiAxI16psSmICxtmGwolyy3gB3VOX35WIlmmLGdMK0lHg8clLymcu9A2Dnn
Mg4pgJTMS3UcMLDycfxjZ//El8kJbf/dYAOMh/2HC6DYJYGqhjSwnIbxRYtKy9qkqEREqyA3C5J4
FTnsqnDAISeXlozq2xvWZQpfamXFHHcsy9RcBGBKIuIAPUcY4/aP/e+DH5e2jhjpykcCBXzqvKH7
p8AbrSnvbk6hJ7VHX9nw5h8os0V6fJvUQ2FoRHTf7gSZNRlSggtt0SwiNrwEC7C4F9jxKB8uHhVe
pAIR5utK19ZZk0CdA95zjyRlgBKJas3k+MWSOPgboZQgBGPrHixvUVNbn/PAxC/Uwvdhhm/iLMx/
wknZxT9wCyk0EiGByOcR0NJazPvkpSrQMTUCi3STXdc3djmLUoBQ52/cpzSIKxJpOROcYDGSMFnA
KgDGlJ75wsX7sApMGBhCnGxnPTe5bvfqmDhsL3N9qzLgt5Bo8ZdR9nmtOa7hVCjNHU86fyrVX5uQ
AqkLZf+qzmRQJ6FwNeZcMYBkJ3qXioYxI+vdgFyfepJLOnVzPOUprl5sI7+xd5lLVVO4Yr6UTr3+
8njiTuEp/1wb9KemTHQDXcTefP5GUNjylEQe3/jII1ABG982v4Stl9CsZtKIHfIVn/mEYH2dEJpv
3M4h+LmTeEeGgVOt9+dbHayWi9UpoSllZrhzkEN3UmNrtXM/Amrhq9DUV8TDaCbD9++bZiLwQw4A
f0Ks+8WdjaxQZgR05JUoNXc9n01lGTsd64knwFE6o6M4UtRx2zo4V+jVsjgb83OrvymzqDcrfmzo
yAAJlwlqCZLo6I8Tq/r6n1pTty7S1MGMUEpeHwpDCsPtLf4tAz4C03YJsdSbqEYrclpImkvDOmpT
J+0bz3NWQBjj78tUuhp1OhTyZ4LHWQiLEMIOIjA6mDpensSzHE7jq+A+14obj1vPFqyu4glbz8XB
IrYIug0MbtS4jVS6vSNm+vs/IMYKe0t7jowqz0xDyLxqTgM2NU5cr74uidut5oTwIyhnr5sGCauU
APy89NSntrMZ49NYPHqk/ii9cBaDWtBwXVUFawOVZs9AaTsCE95aO3JpFteBdKaCjwStCIvKPvLN
m2vk1ICR3D94f7iAt6jvuUplPH+SKJ+uv4sQolKrw6kOLW1ER+aCkjj55yq2L7bxhUAjkmClxWyw
YZomH40Ef5i6tSd3wwtJKXs1KIOspOC+Q3Yt95vKFCFay0YyOBgN1X/DaAEc+R1OMV4/RacoFMbV
jLxpkogGr5u7IY7JGUw66/VxuVtM67TI6AOLDXE9IbWtoPdFQT/dym80s/pSzwvflbuZ9THyp128
78Z7/hIdH7dw+yfTrPjoebHa5J5WSZHz6tT2kduLr/byD01pHStb+/L+4UgPx20Wj/GZKVQzepGE
GyCjDU9RfclkA9w1DeJ/XFnlnf0h98kaugYANmNXDiNdU4v7pJTMpiNy8/BntEA/P2nj+nMDyN+r
bKmoTYhMbwrwmT5ZosX0ZSUH1stZfV8uwyoY+GHtT1LxXraRXYt1TwryW+1RCmv34/AIy9/tRCMg
e9IVGHBJLfYxamqvjRHyqVbp6geWjPfh+JijVUEL2mgr5rwCtxlXi5aKEaOSMX3deD8Y+ytmxAY/
q15fyEm2CThK8sZQ5D3sltssY2aFoVWdfzUAe4cwsy0Vsa9gXLH7DrvUbicWL9KPF9b2IVQro+nj
Enygx5VdUYMwHLaWB/Xn4eZw4vn7sBjknMgfZISk65Bp5QwXVAZZ6W9th7CLJMrnyUG+ohlMTC0g
4bxGAFXPtVYF/6o4DdENYGGTYxvk5iZ8xZv+ubXlDebmE8jthUV+cQ2jOrqg9nd7kRtWZHMmCoe8
GEeQuxxkXeVAfPI2qa/T7xjMfPXWRrJ+1yZjognGyNJRX9V1Zj2oz1uTxM+VA1mTMWa3TtZ3ZVlJ
mq7qeDfRIEMM6WoRmIp3kAGhO1gLAvFGssqzUe4HCVKxaFVrWe0aHftt73fOsN/WBp2Bf+tmy17Q
6FXUaCPw04+z1mg3znH+TprwG1LuWE9eblUmlAUZLb1h2LPljtKD7Pne1CAnoqjB5ulJ/3bSDw1h
KVzzMOL7CnOooOC/XnI0Uh4WLOQpdV2/aGaE/dM+PKeqwgCyG3cbjxy5EIPG7kjo567/T6nwfWlv
QTToIQgvm2TaqtZj4xBOGZF9cjzzz048uw12SdESdcTU77X9n8V9Pb4DKWv1xpYN1Z/9Ok10DyzP
KSV9TTrk3P2gwQcdqXTAEVO9h3suIU3AJJ1I+Q5ISY77VVUb0MxtaRlY9dVUndzHS/RARBtRwBrX
HL49y1r66Eo9SvUTJSODvOOUxxtyjEbB0Ex+0mtuxDtX7Jeml0w4ED2wXbUxUtHF8T5FetHQHbDs
P5XV6vQA0itIx3xdVsFRR+RcM9IPpmbGsgIbLD2w6sQet9etIBWBCXkWX2O9FMUtK4HxwhgNI5mK
1+n/V/mKeB1o+Z7ZtjqpMKktNVn2h+3f3drEW9V5mun9svfL1Bnkob+Z3D+daMugBDBWdE/ue4uP
FvoO6o+uI3ZHis0wjCs1q8jLvdfqv6erMIhhlCvavQEyuAONsgZTm1dir9JfQP9XQHU5uKOxPvtp
HvNMl1CGc9QsBWd6AP56hIR++dKsWYduB4cA6JxF+xSf5CsHIYXq7mgmXI1h80k1JXfdhISrIrzm
owRlI1c8YQ1bXkaNYz9Ws+3f2xkgwg9i1iXIr/V2Ky6Uv8ta2nnjoVUw2d2S0UO5iXaFNF+6wGwc
N4Uoq/PdLY9KxruAY4Ts4e81HKgGNG5+tpb/omBGqDL/xVgginxGRVWTIdpQS1RnGfsbVCZZcSKY
qBUWjVGWOm3kHgKPpdOYCBpBVSjLxUvWHDQRsW6Q9rn6jGkCrpR9PcGkAg82FUWlPNdkAA+aBw6A
xVBb/A817+i8SuXAI4yPBu5p8qz+MdYQUXLMqvTVporNWGuF+bx36lRjdl7NAa2z1crufSe3xiQP
M5W5sDrrfgegH57Pq0WsVIIYLY9zaKa9VnHIQNp4+yCSTlLi/576BiESs9/1lzgPPIGkXoNat0b/
T9mKQ+ep2Unrpda5ZqUH6MJHBxPyuAxVd/tdcXbziDJlOtUXVcCzc/s9DBlsXH1jtiD9Gw4SJrKw
cc90SBlJrCvJmvoCXEBIouT4dDF0Ms+wVqhU5+hpvs7DbsuojA5AT/BD0EyajuSMDp6ZE7siOVK2
kFCaLZkGVHIsPN6r0lFDzklqAIUI2OPzHlPlD2ki4yVNZxKmyV0m6j3mf5CfYszd7DNBowvkdMHW
iyJaErIE5+53c9azB7iAHOeoHt3MmUt+3aX67w10PRDR0nUFGKczE/SNqxJGbA0c0f379YdT7+ck
pOaTPPNeyaRKh8BEQbrkV2uRcmTZ0LdppCahhFySdhsCT16Uwjg5r85lYdRgi9aJFnBHGAt5nTb5
c9zAt7rqB0GRMxaaelh8nfgBbJUPk0Tzs2FowkDOnvnynrXUOQrd7FPLnP1BbkUORhoqqcSC/J+w
Rc3UxllZ9I8DPqo3k979dYfDIJalVHKkETTlIucUKojAc2/WAP/JM/WkHqNW7LBFh8JnPQal+uhr
s4q7vMa3DsTlmJAezkGckgD8AuCuIeRrfzmHAlDn6HSDNdsQ0YnblWryVD4lPx8M+sb2TRTUEc/J
xdKR/+OXntmA4h+W4Tm5oAhEKNgcHqRuQmelhsW5I7rzxp+zPDyG5U9OkOcBz/VeBM4M3gv4Hdmr
wZva3Huq+hoHQ7dsxkNWjaCGqw1TphOevD9oEvUblnLZwcXMDxrhmfyp4K/h7FqhzEsfe+0lkWI4
wKLDGsV6ULJ5tWNwI6oc50vfsJg7R6jHdXapIf4gUDgiwg+s2s5K9WMkffuWdDYWzbJhbk6o6Uqc
JJUGupUj/Pb4eMQedAB4OZyX/Wy2G8UNlodfK5IJ/LGxkEBPZfwbsStoL9TZK4pgQVVuM313fK1Y
QkAiOGbn+QRVfO6QBaXbDqGjYUh4/HCqbZB7cKa1riFSVI/RB8EaGUffv/HW+WjVTtpOMrZqI8EZ
T2PfbK9NB9vyu7W5QHUAXscgt9eRPOZUtW2BLpNV29HubnUNG4Wvbod3VCLvINTfrh24e1NxWLxF
/QpYWwE2sTQkxnMLqlYHfAa1kwxtg6LpbtrptE7AgV15a/C7uBcJ5s13RHJLLKvjJzBy7tuHZ9X/
uh+zuFEmYUDtJNGslALa9F5ll/phjyq3cSJnz845RiVxps8u/GMRTjRqEdKAgMQls0NzXn3vCpRC
QpDNOwOtPVFBYGHLSn7yvQeYq3N6QNAA6m/ZPJ/F23O3pLfXtKkJ+/yt0bxTzay26EEF1+sgrSzl
ggOGwzcarM39K5H8giDhMtH6abYBchW46lUMSswgC+0JhPtCOEXymgmTKDuYoFhh8F35xOSD0fJV
oJvLrN1jvHBHGaTUnlEEOEKICIoPt4P4xaiP/E+RLA7W4+LPO3lhoIx/8afWUDR0GAuERHaoBtSx
P0DqYu9zVkmH2vuFO5gSDB8xjx3IZYYMUVEP4qlIvPPqi12ecTuQ+bwQmn84tp3xwaYDbyYDBF/5
cI2875MpvgDovpb31o4jVtum2GLDxGfyAi5lN7jvnJOMSl4zGsRIcmovgqtfSsrDJoD8M2nxI1M+
aX/SruDAPWDtC2kEMU9vZLTY11R31SNuTPXkj4iw0m0+BZoCvtbHBoTSiHgdG8PNPiDKveMreod9
qW3QBQXeq+ngN4+5svDcOb/X8ooGtWQS8x+MueDbaC5Z5DgqXBHjUoQuKUNb/lDABubAVsOqV7HB
/jDhR3r2+ZlIdfEvsa+M8LK8krUdK/fwOGrxVbHyI6Kt/7tJwdcitZvNQ5E/pZ1gujX21JD79dSa
Cd2CRfXH7Tuz6bGOdrgZUduumfHQfp5rnX+wtLvSjQnMQCHqfbZKq08Ivigaug776UoYoNe6CyF4
UpdZYCseSra/ibiOYbDAI7TjJ/HoZcYebXNU7vVU6+w6baxA/c6b++GvwWMbmM9g2nmsfrWY9Qra
wfRJ8xghOlZTgYTSTZAe9g465Vx212uRkVBgHsmKRVBREnJn80a3vtZtoiSQSJXdhcqTUQa6T8m6
1Caen8Acr54FkDhJ3qQ7tjQSOAF7XnlheBs5UEcWy0lvYnbVlNADPpXHAUP33XpZmMf3Runxi5cw
SMiViwQ23hzba1eUgTEWEFHucMol0MJKjZH7sjNdbTGNX3bcy8gOwUzgq8UdNWblYvt4E7iz5/eS
zWfc++D9Q87eFLS9jHPlVNG2nU24lf8ed76yCwsnan8SPhNnU/0YYD/NCK0nvZ/zMYUxqt0mTCjo
Utw3AwAaZOwx0tUj0NVtCDhjwguEdWfdv04SnEnRJbmbgjSegSEMEoyZRfx6NIuOILF/ZcOd3jsl
5IWcJzCYx1/MHcZgrsB92vBEAiEJzmKVihWUVa2h6IKywoWbZgXElqy1cSmGjJq3RbdNcot1FOrr
GsFUEAJLl1Go77h/I9A9lmPW8rH6Vvnzg1YnstQb9RGoeSWSSE6ItPm894Ve4sw1GghZ7+nR6hTR
vrDRPKucDIvSjWNacF3PKRVlTUQRvtmUESzVYcCKaId1mbfSMFOJri3DQeL68AC3SZUtvYc1biop
zM9vzmMJnzvuvwjuTuKKnHTZwGKlZiGFMvYEtVJrBnQz9DzlSjmy6KuioRnA5+oTppnQEgeRYA+U
dJzSjE60p7WQ5eKiyVljdDnhk5w4QgzcUmaTW1ERD5EN3C8mf+lsGNEqZXuDm/vw8RNRYEu9Q8/n
4JPcPADqB1SQlLBsI5RIL02UJxIKHlhY811K5QFc+dSbuF68Z8tZ9r+5DuP2Ht26Erv+5utBAERV
saQgOoPthTGHUSJyTNj+qp2jJ0KvE5NzRvm4UpdQcbMWMj1IZtNOmiwTQnBCMuOjYGffi3mSYC/b
oeCVo5BcuaG45HKoOWaPN2P2zXxRhMti3avxUdm2R0ZVsAnacvB4eGfoi40tJPTHBljm/9iZ/KvW
a9r+wWzT+P4WTAlu9NCAgcAIWT6VdIQddsYO7f66/5ezAdhOcBpeRrOOjn3CIOL8wX/16OtzpW8/
o7MNzxZ39tzd67Gep9LTQrrYSidxzNo4Ri1/hOns6icYct5HAL+O45LU9mNt6cIscIz9ZvyEx9Mj
OwwuPN8xbww5txzukCOnqOFu0L1mGxNTHPmdgNkXFrXN9ITU2ItDAMOEAxhZL1011LUdwThUt40t
9rfsQ/VJdNQwmqffZPHMsrubfiPgo0omcT+NBKeTFYo2tcdedimpprBOlGjyAOjNM9ftURvo+ZKU
vUzsGXC9eKlGR1fmKrtmGu9zxIwFiMMyOY2Yj6mAEq+rre3bKZlLEjEJsdJy8loTnLwazvPB+ztv
feGyl5G4glxDTCAK/B2fGmVRUs82WYtZpCcFpk1eKI0d0d1xeyo/3orZu1pq+Yzu+EcHgB8gEtPU
DCY3Ng+X70XFkJ5wShK/q1ZZhklW0tefLrxd7pJtMMQ+Czmik1ATBx15nBMGdPbGTNQHIEWxTHOj
+j8N/pUwW/wgd+X0R9XnPm5kfqFTWX4vNAKSqZYfskDG43VKtkxPmMCxRJLrJw+OQdytsW3ewnZu
kuLx/Ol5jjhR+gsXVEJ5L1zqn1qH8cuLpHBVnLPlgaE//ZqioMA2HAzRJPh6bRm+H1B4uQ03xUbQ
X5GjXESccVzNaRO458z7vtZ/KPvQAiod+uJh8Z+aoStG2giTRBYnVYOr+64w1w3X879Q7P/SvgRb
cTinpVRe5KYIRrE5ReGBQXxFie3XKmbwXUPAFv5GMBJFdEjqcg0yJ3uhDKjEjeei4vYSYqW2qrq/
3GFpPN3n40POm5xGMO+uJ/Mek3pIY4JDuC/RfUDeXJGzBee/a9hfoIhlOCQML3KaVAtxx0Q+oiqs
homXuKfnTiFM9uUYDinviM1zTKeRnblITLGYv2o6h7EMckzNo9NHCsfGCPvPvv8ABAMbI1hESU7L
lWCc8LPYCDAjBMMXNx29hQY00JO1w/mseAPQ9bNETip4MGJII/SrxWBOmj+y/+S2rngBDH6qdubd
PH+ansSII92zruO+4qnWsnZiA+46+75ehpKpwXp4h4tJIYuhTMwEOp32hmtLRWTqQtsZoi04Y3Wx
YDocrNTjJVnFhrx6wWxJ7PKdMqlKIYJPo9fx6/THnYPo0iWSkkZqp1Q8twDa3WyIdyLJECbl0oDD
mqxwKSQkZX4WMKXAyda0RDvE8k7BVUB1td1TA1uEyRDWRxjn3cgmKQzC66w2GLx8Km+UdxaVwsQT
OBE8Qz83/cQiiQRLU5Vl9eC3awAeteR5xGNqHqSXBdH48yTYDmHbbZriJiJTe+IGxgvaObdjxmY7
zW3bo4ZdP/C99gSdfwwHTLKY8+EC804jimbg+X/r/DqGd+Z0IihW0T24X+T8eHZBUNXmSPKUIIFI
FyuP94bGuzWTM+WXIl2ythSDRK/5Vtd8S2bPgdFHa0Wm3USdGb6wUMaYNC8f8JnuV+AX+OjlO3Qf
SG6S0r7zEw5UEfEBDBajf8yUC532FLbQsUdl8u1MneDe+sLjZdkugxNpeKpgtKwEXLbpNGALu1Ua
cJI3C0UgaXaXEr7F28rqDxHE0AfjUwwAmtULr3mF2RMTgKwVZbLL/S7PUeLoPDHK11mDR3yXdwdj
Ff8R0bVOpJhIyDQA05OmZp198cjlnfvOe4U46oa/W8M1qoTFtaRcGldRoJhHPq41016fOtgdPiPj
YKLmTnySpzk0cR1LZfxlHhfbv1cDXOnPtp/3EL+lKy7a7aSKU3hSEP1JiWI8Xxzed1UHy2EvUnN5
MRDsBBU20ZxEEUvqWqYqh02WOMIyb4aKkuFTGwGuE4dZU33ziDJqnBJ6tNXk74SIg6HBNbt0YJ2I
aowgzJSMoYx73bIIEFZLEZ3ymXTJz4AEvM0WhPgetqampUL8Neltw+k1CI1J35P6pTInhLOoMR75
2YCPASoFdssmhSZqzqMAGdMqQyAigRXt4qmp1ZEbgleysC7Ybmnmx87r1bCIWlao5x6trJhGoMmF
UO95WOWFh1VFt6fcEBgfhblLI5s9ZwpXC8QtqFWzXW7myMwm8FdwVK620VcMhq9xqi/aaoPCYryJ
abdZF+Bxo+B0FDU9ny9f9miTvtgeBVNTQUlv1vWfTZ3beknVOxEsUooYGM28LTW3oBvbpJcJYhqc
CCR92/m5FcHCg07Kl6696heEqZKU3w8Y9rAnQlG06LKPIYDDgtqo3g96aaw/K5eoQ4lpjYYW/wbO
r6yxlJ6PpXb9SK0STncf5U6rL2PtCHrnL7ng1DufUr7kwandbesUKgZGZks5EwuOb6IP2UKjcPnw
eitYXwbc9T3WllNxDfiWszuk/uow77iiSwnBLIJulTlE5AlAJpDx3yQN39OH/HHLGzw+IdBsas79
ROinSpgc6LiMUJDWV0LO66PN/imC9i69C0zp4ZrHvgCeLDWZIiokQn6H3UMxBnRpMqmuotRblRur
0pHwWV/ZMBdAFFg25PyomZDyNZIsuOGpz9GyluxrTG1GUTX47DPHBzj1378tE409FvQy9ECxaCNP
9RMaD0Wr0u9pIN7PsgJD4MMHFvt0dfIlfgMmh7wgjhhG6quMhCCMSwquNpoNq81VOwTDLDHggJ/V
inDWm9iPyORVIDorwz+S95L1w0APaFoPc0kQKJTxtpQvOezYYu7DhqU+iL3M/Gg32IOTQqY9rWXF
WZPOL6KdUmxAAYh0G3SxfxZAVpP/GeVFyNvBr/8jN+VuYOOKIoFKY/6d6x/Vk9KaxCEUIaLxIeZh
00V46XuOChMGAyDWOerI8bkjzYFhIexKm14djRzK3GF9pPadfCGFA10TrZ3phFhkiqA0QHnV4FGq
ZsBwwpv1UDJV1YY4U2J195z5TtkTmeWKLm7d+oTCEcf/TAarX3eyyClAk4zTAuIXyzxpQ91ZoFyb
QATBnMGosrEFAUHqafSuKYDX2PxeEoMnVYpuFaMmyaaV+4Omzb5l5THsBFSqQZ096KIDPyaoYGEF
Fta4xfPwHqkLCDqH1Efq18rm5wEb5YfXgUVLOh0YpzuYIyABWK2frIP2a7VUksHCoQRZaT4+tFat
DTWqsgcdcaDvl4Vwy7Xo2tF6zj501HAPVwOB+S/zbXQeOsAEhTmzDIhsBBFW/PAZxK9QBWrZQUb5
xnavey+TBYyALs7PQ2v9Vv3v42UGt00efVeAke3zHvqgOIyIQyG2iIAZ1P0eKtlJQU80Rwm8RcAe
bMnjqJU8tfsM7vEncQZKvku8MhCsh+5bHRQjWaV/Wl+YQC/R6HT9aoz0nRYH2G4bhQTrLvSCSizf
Rzd4fx/pGRs1A/6H8kUna3NLcyUiOXVjVpE3BDv0GJGslWUNivdMPgyRzephdJL+vvjEAP32oxuw
KvVlvVlAV9q8uVFRR5QPfcPShIKt8C4r3KVtHR9Esh4KAQro/5xGYzL7T31g353XGDkdKlt6ra/2
vg7TFD1C+4SUqCMU4MjXgRu2H6i41/bYHv4CULiPg+humX05vQLEwd2Bfc2uX4179pju/a2VsB/e
mJN3YZUKiwJ+SuB8imQjzPkRQINujmZliXcSXFcYfH94U5BOrOmxtEXgrLx8QjcKKL9IBOFgUCRA
gTc2M3oODLEuzY3+mpINuwOmGmMBd+dc4kM902bSueayrR6x1kut3XUbmX5amNpQsVGkJJkf/OTq
fVfNTNV63y5JwqeRjk8coS9IueTxymSRKw+Qvq+yH4gaBb3/cxfruQUKANFG6UFXTZZ01CZrJtHx
tfnKaMP4WNkeM4G4LR/+S/R6SY2NPD/HPE+/eXGQ0/yQy5uauBQvnq3b94j8eYtCRcTrWz/G87op
79zXlGhPJ2Diz6+BOH+rZ7vz1SrAbQ1r3kmloBCCqxE80gQKxuJxoDqfwIunwJHCx5Puh3kST1N0
0N/O0Ig6e05a20Ya7SVemJpONaa8i/nNByuE5477fdDhpP0y/x+WaJKUrkHQlzmYO0LK1BMbxjPA
i8skTNFgpv/riGVwwWiR5x2yfADDctiLzpWgZwioZGoI8p82o9r3aHOvmdCQwywzAhrY5rGhntTJ
IxeYKw9loLXrU629F+VicacJ3/7Huvoqo/lcK8ZzqzLpb0HPmFiDvC8nfCFRvc0Vru4DDPf/E1Gi
hr6aimAEylSxZm24iCuqRDzet1WTCRc1yNzWVXSrL9hztTS1/3QEM6iKZi3JkJEu1cYdOiEKQbg8
by6Sj1Md8FiRK1Ho7EUtuYzR92v2yyd/1hSQdds/ls7LgLmnMeXePsgog0gMvonkkJWcZVoBFhfH
vRUlxo5wRq4upmi88xC4+CLDOmFtW1mjVXSi/wd7HuIeuL53eDn7E5Vw/iK2E991xgn+mZu32YS1
E2vwP8G4n16nUfp6qo/j+zIHNSPoGJeEpPwnk4qopBGDkcQxbgfyVkuQL1I8DJ3o65L1FOz+eGPT
+Jqe4/9vEfQ2epQqQIHSkN5YQ+BE6BqjCTOoKtjqnLy9pl75il3PT8IvozxSS/UJ3pZI0YG3vq77
RN/BtJLcrdwmHMDVCiuzSIGLM4SGz+qYLmEXQbsmSlUQkWjRqeJM7IKwXDaQ8OSR5hF+BnhmRRDK
DWfHNQpnAq0oPWgrgM3084+YKAbH6gaBCKqDWvBmfoTuPaAFxc3nDN5h9bjmWBS9A0qK3aBykiz3
5Is1mc7ihAzqQnZnfQ/FbC8cl3w/mpVMeDwrB+OKSJ0LYaPznUJX+PgdlPg01Z+FJpgEiPuFemyr
0yp8/ixZ7uwSbRS2ezUeEFZ5XpsIr0DR+2RSwI7+dr7L2aOnGqaqhq4vSaN6ziYYpALC8J09S2t3
MulKlBp+tNVcth7nALXaFmAscNDuD6oANEGnC+gZwE0/INu06d10IiYmFzutGPDvpMce19w1qUQO
GfIJ3ct1xoNSPGg7ZGiuANS0zpZv1SnBOEipfdSiPsNraKDYCte8XHa4NgLr9UclBc/hY/plOJ3w
BbfMzmb+voJBzbBET1S/UYt9Di3/swv2fyzQbzC5RBg8zN4glg49ZIF+kc/xydnmPe7wfwFKYRfN
tgEPcxgpa1h1FPnyZcg+ERRa/syZnBKkCZ56Y1KVrOtQ0rRnS4cHetOFEAqeA6dHcqO0BA4aNg+2
Nh8HWXz4Pf2ozgvDd179sVgMpOCdvDBBU1EpzMbdJt3ySM6vaZ1toZmNRouLuQlOiMYgAxWXqAWe
MfRHo3IDD/PxrDXDe4pOfLitIsr61gDMvX1sx7GB83sTBVLLpa1BZh0A5Hcn6RLwVpzAwWv9NYjz
kVoB3FCSo3zWo0IYqwCQEVPPTfRyKkcL0BjaKfZU8NGzGUXPNgSLbv5iIb7Cu+zzzEeP7WYqDVTT
hsk/SwkxldDcDo3CMXPGMx5McOpQXY4liaS/xLx7nGWF0ETGAAVHGST+tXyJUvmo2azoopMKtiXX
8dWV3Poy4t3JwaoCwtP/Pcvu+IjG4ZZADTOKBvA0L0gElrGaUiLnOn14+Efo80Ux17tZVlKIxylb
wzw4OlcKm97eovaelJ4VzxwdbJLH/Jslpn/rNhq/z4lgyWTCedWw4fK0jXXFYtf6E5MalVVDP9VS
bHw0kZSgPRIziO0/0cOtSHyIxUWwaJxgWMW/IOAInBaXRRHuBBRcwJX/tzVDRNfrXAAyeYVw5YOE
xJl6c14BlvTIY7OHd6iAGrgvXzmE2qIRJf0o5aCyo/DxgsQISsxxj8mWLh3C96QQJ7RqVlV1FQdg
8lz6cfjLcA6w9pen9g2HCS1T+qBoMixSao2Y04EFXrl3epXfhGY1+vspoXEIVsz9rsQt7akJHwSr
slJgFob9/57TR0vHfoC7iWHRHLyt6WbiG5QRwjyYPCuetk8dWitjw8Zje7cfoY53v/BqOz2QsGLF
pvM04lgbmK/9TiQqRSTr0XiD/qH1YbCYJlc7yyKnZaBf21llV76+9rw4zyfFbhUWJMPtXX1U+HPS
cQvm13Q7yR4Inr4b/LSxrgFimPwgxyOfzs5e73+yBtEpoopCGnUEBZCle3h/4OuacbktKJvFy942
ZOHMf9hNkiOyb4YsNLyQe2MdF2cwbM6Hwb8hBKTxISkUhqO9PTldZ9vhnzLBGSjYe31pRAqFRtwA
4PZ33/Fr7tu1AuZ2uNb/FsRVgzgq3q3oLcuat+O53dpmxO2Y9Rkb0Edb0idcbqKYL5yDLALswNYo
ByKnPrhRK/5pg6YlmaTd314Hkk2MiHgzR34ZouctU4POEFWAL9QBfrh+LfvEQe3V4R0x0k5eZSAu
LfMlk/3xcT2kOG9p1L4nUmKHznbYnBlvuTwfH5ZYDfEDHg7dY3nkQO7sZq6tNmNboQoGELSMhmVA
ye0/IHwJj76Y6b54tQrf6Jgkm6UNUD+7r/27HaPMUfVVdDNowmE+9b4AV8tsV7WDBrdBZpp4di7q
jN+nvqquClh14UC8D/YOZKCromfnF1EeTwdBIV6HEzT+jAEVqHtw0nH2VpVB/Q2Dn1lxyk7g38A8
rLInLNUhxjcqUtWQFeqKia7rxgEzk6YPpjA7N5qFP+vWiRazeqRtu8hUQV5ts1J6mtX4Wsk1nMQ0
RNw24PIAQg+N1FaBOpO0/8GpYEwjz283aXHeU+a7OR4aj6y+QFeaw2p6AVg/2lg9zBLpske78yWH
0UsMHloJAnN3u51CDOPcJfFc+ABjE38x0hkvLgNYBAK/hJ/KWqUnCOMmg5iLs01ZHYTAKfPt6btq
I4EXydtbwxLKIVpo1GJau4m7HYVc4P+fPt8KSRMyvmlqhZqSRiYnDzPqj4m+CVRWLpUtl8pNEorA
uG42Gk7ajtcbQIynm3spwilsXvFrdhQylsVz9TKzPJVDGIlPYHNr9S1UYg3niZTnGdTcHXAYwm5d
mkqs+gkhyvSBZtKMvrMQJ+B/+8G+MmGDZIrjisjVbWd3GIpuZhc5iaQhwsuI1VXuBicDlHgu3g1g
6K0RENBmR6yAwdFi6vfRgYksMa3V7zf+NQRk3N4VaXPH33tnseqUDKTY7vXwYJV41rRtaEX5wpZy
w2HPZwCkzUOI61T13XPSXWSV13eEh6aCORfoat9K63WCQYoDjAEwRpjw5berefBX6laHTf2SNEnl
zCObN//pknTQgIUPfir3+t/Oc8AC1LGuo/hXA6VpdEG6dBi810EuRcEPRRPcvLl4Pb+bMqFkBBH1
j2jjunYxwlSLpgtFcHupc4BKb9bemmvYCpxz4r3wKXbIy2Z7UQCViiZXHgVqir3NH339R7qpVQSg
nO8HYySVHMqrBLhsUylL2MKpU1B+jJP8z1aUsYJM5Am5XsCrh/xG+b5m10raynCPu4MW5drTwqt5
meJUHeq6hyb4M1q4raUZkP4Nvko0AEuuu6AzF+ip48UuQs3qgKkB5xBU7IFYKwK0xT8xcbo3CeL+
hJfWmLlgd/PBBa//gMu+rigF13iZ6EMN85+mHmDbWg4f6P/17MNeXIgrE80dO9NEFQLJnofYDMdP
tJMgTpJ0ULznlmtpMbmByJyM4TrKWnvi9xrO700Xop+25347MTr3vJuFegkmIlRPGcWusx3qrJaK
KCZ4BzLoZSkF1kW52Q9ePgeA/xkk1xzGYjh1Y5IaotrKQXg2m3JsAflizXrK0Oyj3l7scGuSDwg0
+S6/IoquFNR6AwlJfMiQjGlCZFTGeweXRhQtCXNX5C8RBSVUkSNjaQfm4zBlijPhfOuCmmJQr3EX
YQK3aAiovD7mkuyG0BYTtr5VxfHpRXmKQb/55F0RADlDVZm5NQhEShyP+1lr676Eul5aRNvuffP0
BfUoFpAxveK4VSSMOq6G9E7LUCAGUomRNbcuJZgXmnl+k858ZK4NNPRYs4XVWTvzPGhKKc97Pdc+
pkuTeMvTJP3AuEpn09B3ph/IGpbek04KBJYSI76WKphKy4mXfKuKHb36W5p15MHBDpfTApz9k1lj
/s8nUpGJTDqkERZgZTnFdgNTAUrc7aUabihn64RodCMg65v6ZmEBmqwSS6DtYquTUV+i1JawUBSh
X4IkGBVH5NhdVrmZIoeHHO3l78vzixSQyDrbUN/XmRpqtXE07PqxAAqfWKHz8zJFoe8nTNy5737X
bVu6FIddiatBzENtfWa6pcLiqhzOsRtdX+YTplDOih3CyC0ojR0hMy06ZzLQbwGc1F1G1MkEJbfa
RsX1LCn34AE/JhjxXwvDGzy1ygCKS8mIeQhS5/WvmCwhvcU2E7FMsFK3csk874NvaTgHTPNBLF9b
MfZlSQouUY1IDaWVDzJSk9Sil0Cu5pNpBg+UYJJzcPzNimQ2DiHuNpSTPCrHBZk5QXeueysi341r
+sKBh4ha720P0YVdv9i3A1mKWxLljAMkVBPE/UzIJris8JIjHXdv4yCaSUvTvPYE6gU8Ew2e3ThI
FRDOxCM6xVNPYmwfWMBLBHGYj9Ds+u/WCPMBBte/WtxuXCv7IXlVenV6jJ3U5bcX7sd9Yh+2cmZ4
b5HS92dc1uSttTapqMp+ojpBQv4RE/Aa405Fd1pXZvBcs8Ji3KC1Ce3cj7TjA3Lkj8r1aV75OcVT
MwEkySx9QMdmyaYOJ1btxpggEf03U7HQGvR26qfsOYWlQ6ZaeaOsj+/ZFpaKof+EDKo8uRiMsjCj
sRgviDgdEU3HusLySAGw1UHVsXc4akj9V3uAypaCWEGnAAx+mqTTCT5doQnD4ah+y9jllSwF2ZMm
jTog45jSG8FxOTFia4raZowlL2cpHLW9v2N2SDrBCyiONRC8XXmwOIOzrRBFORmDAvJqhhy/u+KY
U3bpx7vu55SJD3OIr90i0J0dM3CZelExrEnxbwP12+4TCXHTDt2bl/QNmc85m8U5VaXt+839fPqQ
mE1mInuLoS+lBxiwDR9s1Y7NRM1Jh+r/qU+4WKPy066+YUD0Lg8vZyzTckuNIDTbri97JnuNxKCE
gghTXPOBa4cH82o53JRw0T8aBR5+hbyASApF6nQeoATdRIqBBppP0QnzYcH6TzwB4bH0kUWVVWuO
5FObo5HFIKWHZ/QwCLvELayREmweDnscW/Lz3EJegoawAUTtyukrRH6x9d1uXFXDBGSmxF5HfiEt
U8jgDaEGLdDhXenlCauZbdtbgPXhLMaG//pH6+JFwTRE/qV09unyzj/0TXundlFIn87Jnjci9x6n
eI3Q5IzPzBZ7ngqgNUQvgL3mM+0m4rQEvpLmNpnzhEG0wMpN7lS+uE5ZNb7qE0B9RwV+yotmF9YU
9y1oSnHi6y5OMfCRBjF+KyB5JU5HE4RjPtYIGpI9Y/9iIBq2riWLwJd8KWdFeciSLEjpjE1vEM93
ZFDjO8rWnWlu/sfbbfDrWEgp7kvbAJUV9lfjszxPqzo1NPPeRfTIZ0SLAJhXyM4mg5Yy9hHagjBK
r12dvUw1YVsG6CIsLp9iU/kAf3IRGB3giKWvTFEjakjOi/tpb3iQwXQ2y0euvSjJ1eGZ0N7JB48X
zXvV0ZPRGGs+3E1eW5SSUZ6qYqbsAzvjYcIXOvUXa0M+GwYtTw5wF/loHkUkS3X8C0YEmJvfctPV
QPDnOUP+iG1/S3egfhXSdIDpKWi8zuWA4XtnwZq6cEHiSDBriOGm6KyU4Aj8V/1sP3EgZ5Y1iwU+
JWJO3ZF4UbireRxLOah0XOs1wPkUcSxfzHLOI+d5cpTiT7kY1kvk0QCPczBvRIM6Ehmomy7WA+Md
A83LuOSug4+wAoqPd8uN21O+5XmbGS5iWkgqLsrNO3NM4n3u7cM6OpiHu5r0c9D24lsXTMMhVl7q
VKgPZ1ALToDT9hyX9NFtuTm0+VT4jCyXASTQwkcMUhb+B05dTqU8YLFOBqfRSn0kFgVfS/hXiYL2
rY/sHUGN2RRxh5KJlQP7icd61EzD3EcPkB6Sn4O/Ye/oPQ0jKK8NOCsOrH6TUa/6B1V3RqT17Oea
rx70JSNAbFqoJSRF7ottTfeNhOlE9ekK+zCev8TNslx34/hHSYN+BKz1U2sjjU3VOgkb2zLjyomk
x942ATb8LZs0BUxlYfs9UNB7LoeWnkjU7x3XK8ernzpdonzCMK/SZPGIgDxXj0w4E1PQnZ38gj9O
YYcrn7DQ9UXNJVXzchjona5rUHOGVD0sIWKFb5mKOOhH3JI18uhJJ8a6ey1+58DrhY1ciNABivFm
+686NEsUBBgBh8T2Lz+x7MzK6S3skkV8TUzG/PtAMCh4uQd3wfH9GzdFuOTusfnXve6IdVPAaDb4
xEZebwZ3zCh0IztF/Zh8g4J3OzdPtercmCnMp53dAvOEH+aC9cSOWYUQ1b0eBNDhQuvalIYolhW5
s3rJjukBEKmpguVExwe/jfFoBIPyDqsYuadEIKhUX7cr2myw5+8Arv1r13uTueHiWZBKodRC1Mxh
R/wsbKwdUyV910C/ivyoelHz1PIYrf8CaFTuXTX8aLPpF66KDMWl5WEAfsFu1sXX+eQN2YEJB+hW
Ha7BjCzWipi9+uPxgqA4gGicfpKOHx+x0prZbsCzQdIMyG+e/mBopA70SDsEBUw/7qRz1oHi5j4K
O07ZEhekYpyaLD5EE39ysJh3ORK8JqLvzNMuzqbgWnu0IXjvUZMC5zuJfgO+EHYq8rfqv/qYkiUL
0k2ln8/+AZ5ZUxy+cSr1rtgw27iQ19AKOd0GgHRoLS03pRW0LFJX7181mF3r3XaTH2bV0GngaH+c
DkoM2Wf5vcgsZWtlHZKGxURqeOWkkaPjLfwnU7eMrGYXPyHWoLgYKQX0eFs0+ovqeZP2/JJdrjtU
8igVnx36k4p//p2LMZSK/vvDHVp6yERRV5WnojF5EgUMbG9b658lFHh8xMLYTUGJ7B2J+5e7OGq4
/gj2sQxb04uX80yoWqMwxUxSzfyIZ2vtuPwmCrb30XAE9oPNqLJohprJgsrMriH84npuTdNueRLb
ykLgKzyIarN7UmGRgsN3pPW++14GsKigb54iTMH/++ul0xQDmZPCDwOLQPOWaVNVH0+TgGY/Zg11
xSKM+XjZmAVrAarDmtXVE+n8PWyu/1TbU4GYxN0/ImaEIWn6AIRZRNlTlh6rd7sT6jp7UoizvB37
o33iY0Vl5FmQaYbu4AdHUQ3jXF5gYEUHube5J+3eEAX32knixm5cgJCZnfYvD8VKaTNMfh/UQAAA
NxaQf+WbD9hvQMHnPhi33TvN5g2ItJE7TYEE1uNd7EScLzMxLKQXBEwR+DI0c3t+jF1Dapj8nuwQ
kY5rWCN0elNpljK5KaSgmuAcP1DLXXGYloBqyUmdAnRxZIEw9/S1I7s3ECBRqFEn/L+PcXMqvi8V
2i1c9b34PFoVuKO2c6Od4oA0bTboPvpQ/NLCRY9oXLvV1qQs62gzYdON1dE8dFfKT5d0XgoFfL6T
PbT2L3deXYsz5PQPDhE3LxFmOcI9bqbTEV5gIXL3Vl8oB7r7B82ihFe/IaFAzaBUKsioTo7Ezu/h
fd4ngWaXx+lA7q7qU3iEdQzytN9vcQWfdn3xze3kGhyyP4QZaPeK3Lg3YyNdzpSOddqNa0B4eKV5
Os1aS/gZYzuftb7KfaT8l9i179sg384QpyPxGdZQzm3yB/t1DzM6W9Og4vdxWYiPiZJtAom+J+g6
+W/Y6zW0KjlnGTPmBd6JshQK/BbaRrjTtTCfLwT3J5gUTGONDBx16Ic21xX1h3GGDAnfc7Tjdt+I
XQ1ZCjfBbbqN5Y4MTkrcXsq4rfjYZsfNq6NXMs5OaBv8ri67wgl+W8NmyRNnKHyP8YSLfAN6mxHy
9NaDmKZfWDyM5UzgJ5Hk+v9Ho6R3h3oUWfJz0xIFK5wiZqB6mANPL5jjtKppydNxpHktx+7zdKsM
ZdVXa8lpgCdzRLirLHlK5Sg+MVk7tA2CIHwsJvKyFbz/8W9GwqLH+MBPu+lkGvrS08m/sy6gLsyF
brUEz+JvC/01abldqRrqaeFts+/58IllkeOSeRJDqaQTaTjEHc3N+xlXxRm+ieo49laJKB/mBmmk
0xoC5oYyJUZ8xQbCHrGljwJNf659Qd0xZS9KhUuIIwP86vQvNJu36nF8OpDbChI+JBnMjo7yS3h4
0gne4DaErvXPORQstqnnE5VCV++qKYeLzYDhYt1r+hEKxrMvxetKkMEYOgx8udfzUrDILyXO2D89
kSm0DWnimd6d8IY3oCcgrv1lMvN85lebuzaZ19dKd+XWsumWkW16uEmGcVek3gAX1cvnAXfGs+Kp
8d6fwXDlhsXCd1HdTiQHdU0Pumqqb8r5VxdZb6P0gCdUCWOfhWi5yvuiI1Z3X4guFBzLKr2o8cqD
9BIH2fUpDU9lNDh20IWxTSrw/KOMRLO6pBSbw8pSt43bxAwCIt3Y0dibr3XJHeudA7BLGaRUWlRE
oHtoMFPi6LJmSg1kUld8+byQvWPITHJwLpKH7xWJRfG4SBYhK16cqcMJ8WKXIa4xWcyigdpkuqR3
x127clJTgZiDGt1/xY80FPsN+53Z+KCP2fJlrYBs7yzdo6XKRX9YZT1dTimcoeGsil/f3akrEaiC
L+uadu0Ysp02nBdMbf2iCLimpItyjGo8XVvIb4SE6yVRiv0CDBqYWiocZ/6J0nrh1KXWkJlHB/rX
lKdahb33Ha02P9+c4UorGvCg+h+gJOWUTFreEida3BT+jd6N4L2w1+XCRSSRUgBr++JTuNp8r+2+
c/+6WV86IVqZqGsLNDEosgnnCLI/RjLd4IxJvWIb+yk2vG1uc8BN05yGAb3wPQ/1D9UNbQaWzwAm
X5dwedfgMNUMwInuPxfKp5BxNsUJUXUsEPE8I8TsaYfB0DZXbnzFJHSxrTPw/EIyRLjrgwZ58SKD
8mIQpJvI/6BwRlU5dEQiC1juSSWK91puqpTqu032zRAcl4dgofIGHw1wz9PednwZp0PeZ/c6mFgn
gvdZNTRTyNzerNe/JY+986oILI7WZu+wGtAi5WYCdvjGvnxgI1Z+MrJHsP/s5JSMiFe+EnwPPRtu
Beq1mz9CpNQKPOZR5cPKX74Zw0jytj/wsqUALMM92ov8YGDqdw9UTWIUSs4VfKe/LC2xAlGwH2ON
3EYVvIVLTAHdpzNod3ebi4Mo2hZZ7EL68UWhmIDnh8ZMUuZp2E8887vMGVnfxaSb6yhPW3+yLY2x
3aY5CuMJyXdxdG+rF1LZafYhRua6jWQQqUGx0eVAOUeFuyrsjpdetgk24+UvQHPmNUtyWvoHpUhb
pAx4w0unfh2iM0aK513GKFjUDv+Ip0ofJrK3I1pqQGA3V4tV0/KuHsZg2Q76ndwZp9iGg3bF2J4/
csMcfibPe6k4DBLWcjN8+c/3JCRXDW7n0omAT1UzSWJbpQIODFqmNmhOjuZGS+xn5GK3s988wRLW
xYA6taiW3I4XQZGqoWriJVyc47PBbnNrA0XVsld6hWcydH2pFC22lY716vW52ICv+JfxxZpyaorH
FBpqrXQ3TduJLPahzt7rxkGzjhzPX3AjRVJhMD753/O3u12PlxpDc27Jn9tqL97gGTwpmG4rYg0T
BMufHfxhUJCAaI+D2PDnhoCjLifA2pZerGLZeC3vd4zYXShWljbjdSqHA+8qndA6NVv2f3Gr8hzI
SSiL3WdwCXzIoxSbyRr67PGq3OJcwgtLLgCDgoAlCP/FLch7l88W+5Bex/MjERevTmNIKyHEGovl
gRKOGWaWPaxClE483x2p1L2aabG8D32GI27EYVHecHwqZcS4rYEfOvVwfQzEEFGVx1w3jw4ouuxf
2fhbe0M5SSq4AJC+nr3xbgiYbggupBygdGOFruhq7a0W4vrrhe1LO5VnhzEQHvZHzkFHE8FMmYj5
QBU2LLCYGlxclkFMjdGbQhLiDPEujMNU8dYMCaZzXESfVQ7A4jWKF2FMan429gGSMqXw41JkhxlV
Dwae08l3jwO3zepJl4xg+JzvtTBhN6wMWPtXnL8acTWSBBHF6Z6Ot5OALVVEAE+0sPNGTf4OU3Yw
2LAarE4uWMrTfn6KSPRtIioyoGtPfVGIlUskdov1l99lif31yVUPT9Jm4mUAKxgPEfVolE8DO3Lz
xRrA0mbFBXXem/G6RlQVjL8vKkC1d1LpfrsQqXes5e7OE7Ec6sge/o7c8nHZiAL0u/REQf1O7i9m
8XYMIB4q93lV6VR1ILBcTrKnm8dt+p6RZ0uJvHYIkuukVzxfd63eW2utvefZ0uJMImxiVIhADCAX
Ru4Nla8RvchmEguj9u4qFdLDnsNv/IPUU3mS8PKQ7gZ69Y4+t4lF61y5S89o8w9zSJZgzD2dxlLe
j+rUh91ZY53TPvqGrbUz16JokDXQhC0A6MqBVjz47GneCVd1tmshl7qdO3sSfZIcK8f75thKD7A7
w51vEEgXFbpmnbMKhr8MiMyDWKjD4Vtx3s3M+PBPvR6pZNuDQvh/dJrXJUGll7WV+1iZ90ilfxEr
VQ8S8k224VgqNQiOBEtR7Olb753yTZUFij3up7jJFPbAppBGi/6U1YGf3GurxfWuY4Tlhp7rT5qy
dXFNOVYYB29Oxu0sHOMA94dzVk2MMmXN+Zq/ceNC74A6H56LJWdfk4sKjIsRzNScc455UWBDH4Iw
t831p4SvWX0J+931EgqP07C800ROSG1tC2DP98luMCmRnfDpJ9mHkKHeI8pq/U7eHLd+HKbHVwM6
81zdNl+NdEmfSE8CHqw40WrBe/tDPSPm1XaqWzQBLazDoaTMuzHhvpzQwbfauA3XPkdwgJ46X5SS
kPfoW1t2gGmbje9+tG4YtuyOjO4hJyI+rM7iEHvrHCbsH6tRFuU0giP5IsOmPnNKzFcz0rSd1atR
bCYHTJWBn549qHsz1rSQdR2EyWhAn8pbB9akHQLTmyzsd7/+33wbEF89JMOTx52j6ftYOUCYmRaq
ugK7qkghjG4GLrzF0EpvMEU3GnTxvSzhydbv5e/uHYweW4OgZhoAE9BhPhVKYRoo54L8l3PdBCJE
oFXQpq0mIyPPawm1N8/CgWlCZCqvQ95KaVL883g/vqmgXzpNI76/QwfMX4oCNOSyONBqmyyh0cJO
yxvxM+hx4TqeJQ0RpHLSqzLjvKzEP5XYErCPjfAZPPD4DJVt/8/88j31I1py5/JHhdlQL9/fH4qF
rSPJUTVbo8wBM5HpX+FkjoLyoU99npG6HhCf7VcASC8ZyokNc9IQwvTIgoOtCf+yI3W2ALTSXjkR
mEAzHi0o+SeSFIV5lDXZTcFITb9Za/MggHsgzIBzxGsMI97iL6mb7j9XyvkAphlnZfgvybvDjcme
eNIx07UygT4OtMFVvDdBHfSweW9XErpPhaj28SS7Sovgric6j6MD46tIzI5UotZt9ubGFK6zhvQR
zmT2duMnqQCbeHhh3+9zxtFRRB8kvBE5dIKFWT2hzzuV4Z4BYBDokfdent0x2tsW3WciVJS/RLv7
x4Rd8pdHZd3LFRhQUfaQvwd4mlb0eJltWH6bHROgE6iO3A2uYf1W+Ukb39dvpk+U54q+mlBoqsOF
cz7Q90Ik8frclfVs2cjIFTE22gt09wJ9dEtnw7C547+rKv7+4VkaM01b8/jwEAQ1c7DK8Rt2yXx2
X8fBynR0ROdDcGBdAOJ8QrGoPKoD+JEX/j8ISjyjP0svnaE9TL7zCpNVHsuuc3craDM8NsorkSJU
cDHU10P74YCd5xkfB+9oOo1TQ5w1zQ7oKmu+04be+qBv4Rp8WyArxwIsVlsOWrs3HFeLjNWVB2FS
wyjAYZBwlv0lNb8H2QfkDvH4dpwSHBZQScan59Uf1Tfybz2lsVUWMNohkIQq3wiiucgrAcqODcZS
/ikuoQzKh4WkYY8WnElYA6VF029tXHlF+8vZGF/96Wyue3BI6d97xLUGNgyWgvEBPqvf0aFNkVO4
J8SUAUsR5JnV5ZHYZGmCE12tx2CNkgVi5iuKrulu0Yt5LDuK//1oiGnvS4RAH9o1nh+vDh2/WXq6
NSQf2n8BKjKNSm9aQc6JPNb2CKzN98uWh8MaPHQrrXjbfXX1yIViXPS4QKCiAhbCQEHz3iOmvmGM
NBHJ6ZFfYY6vmSG/wp8L6oKKXGZSYwHAZMBSATDQB7Yid4QX+0gd5qSUvVjx3CWoGt1Bz/4DRkbe
52RB4VS+irgUvFFk614riouY/Cl6xebS/Os2a7CEZuA0rDXEfdfKV8iDWjAg77kwotDMf1Agu+vW
YZ5RUFUmwue5q66Mw/ODEnkJeNi+geEotaqRb18XRJkeCt+Nzv8KobyXaadkdxaxdOhPkfkU1cU+
klLzlOTv9iOu+tt6WyUxTLFDO2ViD06zPdfzYBLAG4RXWzQbhh5ivP3K/qVmczYFkloDEod5Jjsm
5IceIJQqlffX8vKld/k0J3Wq9cGT6kbt32T7MtZ+cSueQ2lc4NTwbU/TJUmUWIO7U74UM2xDpDRA
9N1FGOObJ2h1hconvze+zqVWNOISw1KyAcxkVkVjQePfokW8/F1ZI039s3MHRBaoCvG0byljp8tq
5KPS0/VrrZzthmwAWH4yObxYh3XBn3J5991cDXQNCBy0PIeLJ/VQYd46MWMNFeKgbZ013DyCJJGt
t64k03KLGlVJ+v65vBcVvrNgqYvlURwZiFqtS5sOkI8s+yvN4xKU8OtFyeT1ZMP1Mkw2zj98SxTD
B9qDay6k+/O6v7BQela8wxy4zg6uFeFAeq9adzv8aFTp+/sm5EeGHnULa7WrLVD7ojkQWyVr/54q
XPIkUvfVjXMcoV5G4QB25jK60l/F8HPhDSdsEy09FW1mwp7wQyhAnnCIH4t/eJWGhTW1d558N9nq
owRVPCYL4MzL4pT4u6heX6e3BGTgWus1HH0v1n+cdane/4qJ0mLYlPRGU9n/cXc2DsJHlFo24oga
G4uMc/zTZzNaWtpaHYJfapFdR0h4Q0RDK7pDgWA8VdGn+Ckf98RedNQ/RjuUzQV90Mee3H6OKNuc
foHK0eXDKU/rrKslXYEBMx7dEscJp881Kb2h7NPQxHlcqLdd/Y8ebp++QUBa5w9lpBumFPMn6scj
iK8jkdl8e8jVGA4x71XgaZ3OYEjVNJD1luk+XABg9NOcdFh9Am3Li3lbSQqkjkjJLx2f1/Jjzgc3
9u1xqCvJkWf4UGunctDNTU1ZBVXtTr4Fk4NW+5fJk5K1v6q2tnnDtHI2WbIThm42s58aHCxeWtYX
3ubaNErzSTJJPTooWr//HxmDJ0XjivQKaax3YtjwcWlMQf0RYFM9ZWYH4+oPRuR9rmyYxpuWcGdx
ONtXcPrPJdEPR75zRtntSQSSideso3KTPynvrMcxJhq1kNCwqc7b9JsFCuISowoBg05/fWW29ESt
rT4XvicdA+JO8gWDM0muduOhG+/VkYyCtS4JAiLJ5FHK2hWfzihnW2HwBlAmcUyn7KRINr/qNcKX
k98YvdCKS962JdZbRzxC1VaRVy8L3aFTdtkubIwN/Wp2QWmqidYwse2xLg7wGSXtW0ir0iwkwFwS
LlKrUyu+XK1BcRaEfTK6hRb2U+iJSUpC19zPhGOv0MIwxoi0Z9Itu3WnS886KqcVK+iNU9QfYAQS
9u/AB1bvOzZGa6V+CMuYGw5zMIvQQ6Z2GFAvfRROAhG7pZDpvbtTc2cZ4IlF4Y4CIGq8mf1QA1fF
nGRzy3Sa8ic3QRZ9HhqbYXg2WTjVVRw5XNiCsE1bkpEOJX1KNxLJpWQtIl0SP/QSYomdhn5uGOW+
Zvd06LaZ7DDi8ev+HkjlVYrKRAwMomWF16iV3iw1bNZjE4P886a2SZ6OWSWH8KkVatJdeSnmYv56
f4+653XGxjJoOcD46IQW+HHQaAuQerdTCYtYaAkimE0NJzal1GmMdj7/r9trgzgg6biNPzSAAKCs
vXXDG3tZAvHTFIzShB4xZspqrJXSbfanHkGZYz15HhVJfAiNhwUyToG/vx7IQTIK2/Mva0oaibRK
xT9FgTVD6c/xxtCzuIUJfsss9UnRskYnjzQTqGuvQJIDXNtmjUbJS2X5vCaMOVZ08zM8WVrcTVWT
cl40EeTfCzMfvFyoFkVzl8g9ynvuNxOfRH9+W3pZN3iAdORkevNtz75k6u5UYu2AQ2pZd+Z+V9t3
uda8kNouf63tR4FTuULvTiBv25khzQdIaHcF4Q74Xqy/C2vV0Uu3MhNBhJgWEWWuFISb54jCbLMu
pV1krR8YbjB5wAcOsW4qLmhgrG5yvYaURrqEsq+ZXLev1jJnoopHpuA829/o4bQoWV5XspZA+/Ay
37cLWZvQS/PuZlU2rRR8X/xPGQ0Lpq7GpcPVhPc54uznYNM5EkvnTKK0KDhYqKcddg8w5T7Cynud
s8yFOZI+3QXFslfJ87kTdpWv/s0GfK0wLqH9TOvw9rhy+I8nxdgbQMJrHEbN4g0yKgLwMBXW22Uj
t7SXukVd57LrvEGPlss4CAImlLb2LUcl3dM1t/C7x8gT5UfHNI37X9dxJDf1Ex1JU/suaUbOGWia
N3qaUF4jPH9NZwF3T/fszv0wFC8Z9leYabwjLIQgbmIVRzsVoXvJdSux0/aIp8Cfj3e8a6mRMhu0
z8dP1dohk2X/lSH8Xj8tcmy7RQVF1MFAH37NIvGIZQ0RWMLgKuR1xf1wo2N31dYp0MOjtDkY2v7F
yUTTKEoWv7mxDRjrCgaeg4XGLrdGJnIp1xt3XTi3178S41YEXEPfZz86MPsYt17ei3kckUmVEjD5
j9rys2JsGgORbggWmO5LqPAS4+F4w1EW6LQASlvW5nLfu19+SnQns1Etu6+MkD/mT6maxWwkpmMQ
pp1fS7WPhZA8GMdouSByYioBCYS4ZS57aueNwZY1tDF6VdxndHsZmWyw6/dq4SPT3qgwQjz43jPF
PhwBVZfv6wEcinIAv9h9Cmsl2PaMFbkcl+b+nSshhXDOwzQHiD2HaYc0Uxsd5nMiV9lNAqHGflPf
ZuAdqJxis9zAv//n6xarzMq6m2ul7eNjVMWLeZDhw6v5HRAJmu0zCCGGcOb7qL59QPNSlCM/bFbT
M9OcAfFNZQH7X4yQKWTtIIcbaudXPYIJ23mZ7gfPcQL7qtPXMTkCE8d4keMHIauJO4ZK+zbd9bai
R5JiQp1my74AbNuvJKij8v48IXlKRMFeSCIJUO6EEYqDVAoPJewzC7SYqGB/akPTS+ZYZBdSaFnc
fGyPZoSChLb1Owm/Vp0lh5FeWGBqMPSzDpMPL1dTAa0aev5Dg5wGhHogkGRAfLB3tSu+eOuCW07T
fOaSNwKUahmm67XXBM0IOhg5F6uHiuIWC7TkpVI5bGGCQBMF9Z03V0ta6R+OOv5HMbCRxqEN2mb5
jNDP90bl+G13JhkMlnmQag9JCtk+jFBLNxD9rnRkkDdq5R2p+BhOKQsKdrZu869TaLsOSwBR05AU
vNDrgoogXHn4UxD5/prWNfQAxsDHQlz2jzzYLteROS8gQ9ngCL0DKnVdrU6rPfH0UTRC/KwX4r8U
J9EptV0GcYwX8LfzbsOFKVlQZElexuriGSHSxns4mnyooUp0eYiK5ogQ+BqtqegfbF27DUPR7+K/
Kxb2qpb7LstEwQUybPECzmYpiqzu3t6dq+2nXzlF9Q3b0qWxEo5399wRPn5/YRCIoXwds/btgdXa
5W7NdH6EoReqSeGY0eSKVBNhH0Qmc1ZAS0j09f+hj4ZMxBEPPV1vVDDgStbFDkufOvQ2xZqY8sCG
rXHr4cV7F+8Jtguy1Lt5t1m/hDDM4219dtuJcAbpvPZGZa6zTWmdHP4dTxn7B2Elu84k2EzCgFbj
0KdJaalhe5hyzmv5XdXD7Nz+659jywwWGvPmBqKRsmFUomQkOv/ne8Mb2E+C+X/yBBZurs8Mko+a
KF0H9aA3LQ4Npsy4LRZmwX8criRC6XZtBX6kv0RwteACD0/ETMXD056QxvKo/KZSdNkTgn08qGg3
GNWiS8x3ojxDTZ5Nfpkk/unL+CnhtUytjo6xyFd2xcazOX/gUQomLVJVfOVV0qPROgNZ2sqO8Cdy
dvvZoshChnjbFHRA9GhxTOidXHBU5crX2tr8Ns2gceY2iWaEDjBsrEzqcpSDvL9wChBF2zJeBzoQ
zb8q/zIg4u2c2Fqqr2y3Cf23uDiEazaB04cNWmkx6jvRValSnx/T2LyltuinjMPSpw6Rgrg7YHLV
otdYBmabbYacl7gdtRTguIg+eYF4SjjfJhCjJ7rxjD11YEpWD++iK4oZoSysPVsHr59OllxOOFPX
lnl9jAZrybB+vddK2Xggdw0645qhSFxEemVHKZ/4SGbdIbBtE301FVjeZE01b375NR5lwKpwt3Zv
8GSEJWJo+Ehn1uiSn82qSB62t5QQlO1cDSRbnuBqb8bZQw4Upt9lIT3887uNRJbFAOHoCWeTvAn6
I+wGuGtKDrDMifXx7e8oABpXA+9AUYyFss1I2DfjXacYP8+zx2+GnJxZVG87K67iLu6MXG7gpVHj
K0U1urv+7+fiUJAUlkIMw2Ta7ChbbVrUHv99kCppGky07tcB4oWQzOY4gUrF2gb7pM91V70RAOq5
6anZBWAOeDxZa4Q6j+ESHPwPNTIuyQEM0VBubGIvl8l6PM1mfpdGzUg9gV1nkszGHwjCL6dEura1
DGgSdGu4JW19B347GFGBoD3xj/DCXPZrnJPYrdbAqqIO05IIjbi0BjyZlsxtk0PNbqBtOiadTnh5
1ei/cdwN49OyLoRBNhPFXb6mfyQe/rkUePLnkxmuYFH3h2OOPW5zDxqTmg7d8dlRUsljhyPE5rxi
zqJNzNEurrrkwHFuxewL/NMJ3qlX1oozwNd3nFQnvNtgrHmflkRwvWYblGVsEw0zZTw2/fBIgQZ5
yuX+7q6HWaRItam9Nka51e10p69jh5KCo+Mp4YUmKf/MoXatsMSDjG6X/8oLk8OnsKid2QYqbqLX
3xjGdSAtQX9Fjsi7hWj218/MxneN9NK8UQ+aHDS+t3WWS47xtGEBkVLIZYSw/Hys9gw5r6aAUtXL
boumfbUSZxR0hgUz6V/VD9xDkqL9LM7PXQMlet9qlPkc2muQLvWtWPePM59FCk9gR2C62DBsE7gl
Y7swak+rIcIoclWOuvmgL0zIOjDU4PrJyssyZOUwNYURldW4kCIJQIuvRdBWcMH+IEruSFJUMFJw
IUVohhOIvQoNQhKCfD9F53sAzrdABwdbqMEnx5KcZwQxuVDHH1/MULHxUN2o7YCGtgHwa45uQGhc
eOov8YrgtTdZvix7TQmdvN3sFOB9F9lTOpQXrU79G0DtUGJsaUYGuedpXTlH+eM3GebEwJLuHJVZ
MycxNOpgWtDSmWAJfrjeL02sSvevXY2TblZ9sUolKh9/0/CcoR95yGVdbOj+dU1pxQeGj1B9qOhU
7PoL28aL7NfSRUySWcoGaLlWa0MpmNafIjYJy7Tw4qIN8ku2BT94CBmXRx8gWFtiOUsafWiT3ouP
tyImDBIYnmZc2dh3N+onUsY+icoe5iGEShP7otA5dUSXXVnyUUzgsAQIVDlSXCYHzG5/ZkyXsouM
VMK+G13aliZUQjZJ3cuHxwsySMvkr7yew4iu3oKdgWKH+jVTfMS9lTrPP6NQijy83BgSPr3pOIxO
6kdVGyeBaL4dvDjIb3X+RAnPcowrpamo+3GVrnaYCDSLPm/htt1tSbsriu2GtXrm76bZ2aDpvkKz
+Hp16sN49mG358Si0E/mpVXYi8TdGDRWWH4NYtcoNXkfP/JXqXPDFKZeeIiFGDR6mILQlftaW21d
amTvDF+DZN7JlnnaT5wre81wyUlvFz4iLqX7TOeJpWmFz4YyOdw5/O7csEmRc1q21a6Yfax6Pcma
BS3+7aC0NTXKvRouKuh0//Xf0Rf0Xa4SZA3nCgUgffbyfEH7yYqmkb+wvInOtlBdjJH+fW5rF+ee
gRPlOv9cBiUXTtm6Kj013SuaBwBoSC3tdK7Zbpe2gv/S8CJ/pN+bxjCmTVyE6xZdadurE1Xd3MzI
W1RbE+AMGhkmNG0yAe92BHWTfeBXBhD8Q3lZSCdTrcexiZ3Bng1AySZDhm/euF16lg11SjTU20Qt
BJ1t4x+RAWurTp/NY2VQ4JDgfaEuPvoMeqvUE9KGXhfThIDNiIvdYN3i5IWuY2huK097m7Yb7SeF
isOF0SUTkgPmYc9OEIQGHfm/e/tr4HK/Fvx26mlnAcurrE4g1ybOR22Q2TWNZ1KjXZwp+1g6U6zo
fmIigk140UwWJejxR738ON5Xgwbe6hGIjJ3u3padjAwfI3yolq+akfjUWYpPbj9yxMIcws6hQGWu
WVPHWiCogoCNHsDxq+JSZKB54QFjroOluCrraX1AMHR0tTuVuMpbW9R6ZCYPp6/QwVrPUMNFXdwj
Hy2ojHhvBPYesBY2zZoBsDEYt0PDkyTXvs0T1rbxPGgFavcnGYDKMbjqn72vIUv6q/mZqHLjb4Ns
ddkXBivGXstsBZPx7UTq/KEtlxGrjNXtO5LYQKbAZQoZvNdOR6U8zN15j60kZI9MlLHWH2TIetxE
JMUN6RZO+HUt3D/o9KfdT3lU1zVXxNioAOJwzeM/QuIKTBDQdS+w6HmT3gWeTliS98sa+wT1ndI6
lhYBQhoWKe+mcD+AewK+Le9N8TpTmOzVqcLuPtYdNOl3wP045HoJxHEuWRD5gplrbu/AGYMtLd5s
1Vt86CRCqrsmK2L4gCGKdNrn3eoLa6+s/LNTZYymxjxY32KLhcO6T3nCvF6pbWva0ooMqG7jA2D6
ChOoRqOGY98OQF7k8J80SBVEqP5l6DosmiX/em3PDWsWnt4ma9x8pFGJDHhEqwist0ins7dfIL2I
XNoJYGq+UrTZ25v3Oi8vp2U8cphPWhYIzByJ+mcHOp7xidMD0LMMkPvqFVzMOA+MozcCl9/v3QK5
iXWHae/DN+uvBRFQ2aMhLpbLGv/UAWPLTiFc9FMabBH9ZU/xkVcZFXpwUxvTHJYSHo5NXsotT1zq
chv42+4SL5Qi6qG449X1xeZd55mXS6oRQNpPcD9H/xivIpAUCsl19QVq4Wm45CqRGXeL3F5Xkq5V
7bON2t5MsPDuhaNNpqwZnlMjN5olGPLuXgHAdEsMZtzS7HQhlcSQowBBWZTfikzyk+IkudB4WyZb
krq8noxOS1hmNgV/2ozM6JcuBGtrL2l5GkITzp5on0Rt2O9YHIE8I5/0xTY+1VuyNvDd7yNPbRDO
ipGVehlZuNfQLx+3fS6jVoe9zJI7u6prp0Vdqa9YN10t2sJodt7HXLYrme3Sbbkteg/VrwM+z+Mq
PJaveLZbrd6UnNQ6cxSQBpyITaJwAlO+iyMnlrYfsdy07L0s3CCNmozqJZ3ws5oY5ZN2kfSlxCMD
QnY+PZlVcJDxbmeyYMpMDLU4Z9YtnOlmMRkDSIOtv7gYGNTOD3fL9VoWoPuCMbs8IEYXZJPJgvJ/
rlvGCM/bGgNJFOcUZY2jskgzGsXTiCfbxUQlsho4ajOxW7/hkIo/Y4w8QL3rLFVY1YHgYEgm8ioj
S6vjjcO9RRs47LfhoLSB64QT0xbPfAydoRzlxWvkM0a+DvlHexrFGOwLmUCjYjNYvVqaZZ5ZX+KF
E7uiLG7VuAwqOPcoejehHVseNlfvIX8YiOHNSCvAgmapzla3gf9zIBNkIfpnQiYXm7T9v3J11h5P
FxArCNzv3PnPL+hedgACmbpuyCLT1UDe9ilpJuEQN19+xMaz5A35/GgbJQH/n26V+TocrLLIIcwF
evH4AyfQQw19NurZ4PuvBbxf5YMO/zgdj+/c65ghxNK3lPDx4X4ZuwIgKVRqFui9UctUAsx0Oyvq
j4e2jmV0voG8cMcQuT4wNUAqkK1i0Qi04xWW6gAbEFBXaL4VGTGITqSttF8hAbEYCkZ2xhjCQqG+
fciIAppjq4dZN1h11QhDeozDs2/ccyTk+IpJ9IEh2Jc6QlqL088Vo9hyXVH3hATtQtB2MwziMRSD
8JAczfQ3eDbJRO1kDYR+BG/5h56t6XRoF1xBEHOG5Py3ScMFBjqzl7Om5eryoH4zR/8pfu6K+krZ
s/jO0OgGRvjUi1RY/3PFhfYtPdBIjSv4xGUsecM2BgfTPiLA5vg75KkKWdqWH1NJQILFiHoC3bMb
6/36Bj/28tB8jjBP35t56pO2RlUL21c97ZSxjy6Lf6o0zDqd9gzkqA8tKPjOWZEoK9EwwezmlU/E
MT/v/fau/XgvZBYKHGhh0L4i3UVOt4HV0ED4+/2hVgQX+glSXKubrByl2ny/bCaUUZw2c76sMy0D
nG3q9YZ/DEgRdaPgekkQDV35P4NAIB2ipvve6aHu22ayU/JcMbGe07TNY7rdX4fevg397+z2SRAA
oVvcSkX03lWkguj3WIB/CaOvQJZkGOSjJzPJgvlQdttuVno03MLcMxwBwb333amMRAlvXjUhnt3R
JQSN1GKIXgTZQcN50EU4eY+3HMncXwjbJnUK9mNsl5fjh29BEnFVPa9I9EcwW/M3b0vfSkz0Hi/c
O2w9VSSmyVS5+vu+jJezRGATX5h6erfoCu+ix6pQ5w0fkxRLlYwZSbi0mRzLJJFtTr2CH3VSHijO
6K4zpFNvtqVPGTy0zK454CUX88shQeQ9hAaspdZfH5JjAX55iZ+xwYK3XYgpmlEKWnH/RlF8Q1Gx
hAVuyBVq+pnShfddjj3CIeUcZXN2urYK7vbg6XPvmGl9PY875yLHH0XZf2oHkhuZ2p8J/N0EJ6ae
9DByZvI5XNlBH6CiI5TaSbevDKaQGUOMygZ2DebYIGfLSkgUgh65I1ROha9WvW3O1QB6ti64hHu4
iJztcUx3bHBZavDsY5mPViHWonH/9r8xEN+yhQU0tbHZ2p2ZwPQEsdwPHsCecKLekUWCw4OykENg
7JQOwL0SrtzJW2VHdWi1g8/XrNYaA97FpY2jUBEoEQOs8mSWtBtdyRipdot/dEPpYBgqltOr4/RD
TwDrPK7z2yto8zfk/1PgIkyFEt2n8RoOdqP3JyE7oDKLgpgSV9llHn/z1nNzCd7KtoJJadVb14t+
lUtn3K53C4BZJEmDWCVMC13ao3TlaMfLNqu0gtOYsYIeWNOQ+DzJ7PHcDIfv0qKnhdyMqiP2J3kx
J0yN+acv2Y5FFw2fIYLm5KVvJgCnNEeZalwLAMYG3h+PhEn9FXsXLxRP+Fp6yPPYJ/EscXdw1/KE
/FVgcMTOUzhodXBNcWeyHGVeSc7RfXrtuCL+wdwOM4z78bZpLtmYpeOXL31aGXfeAyHcEtscEXyS
i5D2cP/708mQNvMhARz4dTvXx/jhIVzkLQfsxsuXcddgOknyOnnLRBttgxKPQwsIoUD+mu2V/Lm/
0LipdGV08jBMFebNk9kumqHyzw9AM8rvx/UEN21CC2gg2XvcR9Vmf+8P92pzwRRxaDnbJLjeusRE
S5jSk7WTM3sVbS7MlQG0KwioQEd44GmiKJqqJx5UuhfCjyyE8we8i2VEyGbOepeSPfXjuTHiufi4
1vEXT+RVNeyxhwQm/OrUOHbiBtaC9Ed+g9ExddC2C2Ws3YtOS16dU2X6bfCwCxjD0dAgsIfs9s8A
So8I4TYodWkkv8LUUf1Uwd7lrIDy2oxuZymWuu07drEiN/PofXK6KpxIPjbVbHxNzxuZqkQzJz2x
rc7YNum+7o+eIIpM6CNP/KzRKNd9ENh6HT/Bih+j4SpAtZQsZbNimgsrGuo7QYvKvTHSt9SC1YWy
XI16pRWy0r8ukQINtq72g8GK1yloQRQ/2y/d1fhC4anubCcHbUGNMdrbefXrdz8QH59e9Li4KVx5
lubGFv6ZUh5Mz6owBD09bn1ou1REjNuZBbov85Y9uPxApcGKslZVNyzZU4z9EEwfxIeOSXhxzhzo
uqUa5IskTJ3xsQEt0j0Kyqh/zpyB2/7Gap6AH1AhB4owfKjzHuhRp1kKhco5KIarZj2pxUD+yGqe
YnCgcSKZMKID1MfxkP6fBiGU7BBF3bB0kz9fT0Dg0nu8izmb9eh1tvZEujsLZE+iNZvqqDb1mV0Q
4XDwl8HgeAvCHN4s6AvONxVsjTTOOL7MV7A+v7po3e5VuMaRQa+m+vHx1G65RLjmJVO+Tf9AyaUE
hVYmtuB829Z3uHKulQuDioeVvf7R+W0ecfbcZ0Cb7QwJAmX1cAn/O93QeZTDpm0dErXGDW4vIkoB
E0e5/eM97MjFyKe/Aby7X0sAaU+6VcLwuT4nj94YrPCeihIdXYpt+e6ioy3e1DHjeClqopt2ha6X
pkA6nRRGeh4l9bf5ey9qR6qar4s9QT+kptFibz5Bz6upvKVxByCqfLc4cKxNOqFvRr7yGdh3BCbC
EPADbcbu08qxObItnjotbHQ5glVJi9R3BLuDPzuDJ2XjKLGuslPSDyuNefbx+Rv0UtoTQ2yQJKbz
GDNT5DkK3GSmJZC56ukOvZpDXRi9X6GVn7citTEgP9qSnmE3ZBUUPSKTMZOOOlM4t5ZBPsquOf/O
vO/JxG8m/a9MXs3O8VCKhDOBt3Y9pJmQMCe4X4n2woQBtK+rUfLnByVHNcGRaFSafoZpOMnB9dVn
VxUvnKEStDH/MJn7YNf4hT9tbHeoD8CzsEMRY3bFAPX/9yTMjBG0kaVVDFxapr5UmWDk3YSZsjCF
qXUDRMsCxmasjZZjqcGWR9wJA4oagPnn+Eovo/FYXqtRoSA7oHaAYP/nDavvj+DldxPZ8C1p0lCD
dZvgGHlVcWEZ3VNSiOyzL+A1BZUsfZzbQUCHE51dZqi9dwpdciwHJ11vZvJTWZaKQ0Gu7+WLq30p
2hgIJ1ZpIqPbTey+eeqxgnza6XBbwGFP6D7rG6mt2JVHZHSTGbQ5ro3zA5DtdEEluxpaGpmcFFJy
Qg4dLqpHwmuAT5IUzdAi5+V9jdKEzQMVZgy0fLfuNKeUPbDk6JkbaTQANFeMHFg4xKBX2Ne86Ws/
9pLAn/FeZngL6G7e0YQM1op8qmx8lyP62h2fGlRR5Clmh3ywGgCF+NHYDSGxoLxVIoMPVDypQgkZ
509URAm1Q2+VNq0YDXW5YYymdnkL2vrkQGJAH+aSLJDiQ8ezF172xf4bCG5g9cbeSj55METqrYtL
r5EfDlbSAdYUhYCaNnwrJOdycx5j8i/Jwqb2O2A9T59bp683xbeyAxMirDLrf2YGhyCX/sp4eaYu
1/+UEptO2tJARHyYyERlakiketC1euEnuy3SNp9fSqHm3+EoQiB9uHF2huzz2SZVuN9cm4n5IKM1
wkoD1TD3676j2/txzRnGp/l0GBWde/4D/xnjubCkvO9GlfUGh/YNCAQBrVGPpg+sFN5hUOcCgno9
rO0/JjqjwETUcB2aaQf6AAr3ydKL4d2nR4v5phO1AFYYe2nUF3BBGCvRoLJxJpD4gPnqGP0Lqx/m
GZAiwOiABxUGFLCfbS/kacyZNW5QR+lZy7AKWazUJ5/KzGan2ZMd99+i4MRvRfWRYqECDdBsHgau
6jkC7+B4hoVsZX3x1moBjrvBQ0DBYTimCKkMUqyGCti5XXw3fdM5Z5wpUp/OsNT+ktlT4Gu7MKLK
gvjDq028f1Kg7Oc+GIA0EGgFM6T5q4qbboZTi91MXXNjoGD8udEbi4syNshiIW5DcEX9PkGFaKsS
+GJ4r0dCk0KbG6Gp9EipXCFAU20YZay1QfU/nzkkd+HBGYqmWFPvebB1RNN4Pkkczhwl4zP2vnOG
6pkHKeYd0ImQb56Kdcqlm3nSaVzsF2dnt8+2jPlm+LBsPwYwKXy+qixmR7PwMbIezO+jMQS56wZK
flzyMa5r8THOImniA2qbw3p5tpiMlJU0oSaGaX0OocbsHf9BBEnuIm0YbmqJldu5fHoyxX9/tjNM
R9aq4lB75zSJfMIRkELuAxG3TN0OkWk3jGxznabQQ/AGVN4iHFANdmOdbt6lozCkm6UalFf1XZQp
7/pfwCXvYeNIck/T2SOCd4TqMerEYruAWI2xvxxLA335foFQgxE74Q6HdrGD3nPZWVxwMN4HarGX
JFl0j6mSg6UuCDmBpCZihoOrmDDhp7AnREfshISy7SD2RCN5aCIlyhYACq9n7PUwfMU+1HHMfvK4
xTp06cM/kDBuTfghtnCazatPzYTkYFQhq47CFi+Nhayfp0j1c1XK6iGZNhCvi12YmtNfXytDtwzi
R1GPl8JzJboodx7CThWtzLUsE09qDKlLRNkSIpue4fmPNRJr/9pily7miq1ZfvrxmZSb75o4JoVn
dTEX1ilRuqKXJErgmC+5Jvx2GGwLC8wiZYfsvwbFT/Q3gWlUVjrmUkNcnbzu+kWa2HZDzPJ6r+Oo
rNuFHHJZqzjxrh3XiuILT8omMzVOb/LOVew2FS+ErUiR7CrphDpa9+gXtzJkJQiDoW9ifJrLDIm3
k9w5PsLhLM/m8z/Yx5ih/jVBwFjsYZXxdlxqOO/bLtuP9WlbjFCU0VFg5T6wBXBA90bLp7pY5sNL
RpQ+r9VLKuzEE2UK0ReSKyukj618A7NrcHsyNDJFAgD3B9l4weO2K8hu4+TTCQ4QMrmVbHSSjtNU
JKhXop8Qz7EqSQSNjlZWzlPgiOrTz76HR9Z6LIQ6b8B+x8WGdv2TZRH1/4rKS+3S7jF7BhcDDoqh
CXg2ln2oUmrNn9FFjBUGPVkzFoGWFMPaN3e1+TESa4iiFui+ZCi4eLDPxom5bKDXeBJ3EY+nJqYK
aImdSt6iIGgqkjsf2jI6/4m7cLvZdFvmT3iJKRmKbMqq5cka6xwAyGK6p9xxYv/cMpeHXLx+Ptmq
WPIgu8tPrEb8Y3EBWx1HQJ7Zl3gJ7Qc2ZE4V5+sLL+2Cv+Hy+IYhxMzaUs/7Hj+OtSx6ecfQHIqn
frvyDzJF6vQoGzSipmNUpuK5HeS+/HZoS+O2MDXiyU2eux7NPKY+tZsSQS5g1CmtfNxBIM9l9+8B
7zaX9oJ0HzBqjO3b1iZgmxudtcLA1ocE8i3btSuT1p2BAd1hsR54e/cOT97T0eNGfj9iIGePK4t5
OLZ0Sz9U8Uxravd7bAjS1if4lHj95wZTAyh2WpNb/4jMJWZ/ExVZnQ3wqd+kWPlFiL1LBOmknKbk
UTuarIen7GWhCDU6kee+ChNUE3LsO3VIUph3CW3G5CoJhI6Awz9fO7nZhAwMBxnKIqR5XQl0JfTh
awzwRdvyC2dAspm6yZb0dpLIjFzs/uqFEai2cNDvpry4cTJkIBrm6zHLEvPexUYDxVP0x53ADt6a
+5ec8Zf9ZOnkJaKTcXNgjm1oqW+gUwt1LoD4U6MHberq8eqrYul7N0/orqernUDNL3PXTSSziMmN
/P//LHdtDSJYmNSRyapuJPQIhufAfhVAPrBgKKVAG++VS2n1gru70XKQNu2z+BSFaYHBOasMedF7
+COJMXLIOt/Qmmf1rlnIncY1mqCAbfcOflg42Qh24rEpdYEQmVt8dw/g+/x2ieHTQFXVvl58gy+O
lPRijktZPlDe2k67RdLgYEwANDCD+dsnxfX0rGcPdHJS7qg/a4h4SyFDtDVzUjTiXTBnKPp1pesg
f++QY8U8Gyw25ySdWx9Wh6GmXzLym2ly0mxzwXFiNbqXEPoj3kfdOadVFxnU0C6lWQ/nVJ2d7ia9
NPYSubFBntParjm+fnStmfsI9F6HTpdvEmQY1ez8U/lfXmODXP7lOGpeGiHgmz2ltJmzLm0We+Oa
NXX2j7T5/T9akC8R7mSUJh6vihlWQLiaRpAZ54E0q3lg8Of4WLvNPLKAC+OEA31RDj9kwLMZEClK
yUYMrgBKwBTGh50gZ7kIjVZE4QR2Amkx/olpKMlW201Nb7pISv/3mozaVXhQ11wkrwRFkAmBtYr4
WgLX6tzKOjMmeUbSk+TZ+4vkQmxW7/9TjvQ9/16dudEt9cs1dB7stVsuux/AiZjGev72Fj4nNNli
Ma0fhDGyv0lq6ybhdsPYUddmDuoMAIJ80c7r+CK9K2jZYQ5eEydvsHgi3dRnFf0AeOQV4ATqyRu5
T2HlDKnIBNQN3gxkeCRWM281qft1pEu/x3Q5V8EM4sueAx8GRpXdX1nZ8RF0K5xl0Cbf+WnpSTqR
pdhBp8a9ZfvWAu/KKM+Z/D4/WYnZ42gskbIYtokiBRKM3M+z1AD7ZuwXLue9G5ODI0IlOTG3MLF1
mRE2T9R0Kx9haGtMd817/RmXoF2r1fOT6Z3EJET/WMvLZy+iggJOO697fk9m5hp4ta5B6Ys2zkC9
3hSzr4u5CtG2a4AVKrlzsMk1EBwCGegIXRyOVpTQO5oXGeOEYaUVN9WGyq1kEPiDDUJGcHOm9iE1
BH2347NundRsctAZ2pqDpMk7ECLQYAzwXif78ByazXdhH9+RFqd7Jxr2iMC9smVTt2YCefpWkPCn
pI+2+Rpd3PJyDhpHhHYod3jWdC/FOwudJZobgqMo6phxpx4MQnSt5vjDXL4gHk4f0NYuHPAN20vR
y1zMJw8sHV1+YUseVSrT2Em6aLKO6neTzQhOMK6hYYjlt4RQM9qAEeeyo7ItBCQ781pQZwg2mtdB
TQn3ncFyttpqUEDI8j93dni04OuUjkrgXgZSoY3Nv1VKr05oTHci93MwTdh/Hs0tJQgLzyLqfKIn
1ztbTSBBwg5/DNgkBCsO1Xd/2sEdEacWvJO2J7qBJsKj4MiRmv98iujDY3hHO+PYLvGtc9zPZ17j
dD0mcaY99ai48qJ0nUmFv0ghHPRZyDCI13sOTr1wSfetiyVM3T1otedGzXza+okSA+wroog5BNua
6LxJPQq+FhH9mD2xm6yGUxDsvcXZ281rgpDX+hm1jbNR29/RoXj1eOpSfJbbHsFEtJQbnB1z91mB
/ObXP/axaoefkDmSSmm+E68aOOmgAD4aYy/G9PuMcexIlRAWez8mzP3+dx0LVfFn2KGGMuc7C5rE
xHGBEnuOaBGfEQPeKC0F8PNgTVoEBx3PwhOnYuUXoc/k4JNvmZIHrblqcxNQjilO11/epqTg8/PD
hNtJCGCE6E0qU2G8RpkKcLSqGdDg84R4ljE/bkak17SFMxhDPycIVChk+D77/4zX+JLYt56U3sXd
MChlR4D6FixHTspKLDZHsiOhnIY6vD6FFrdDGbbN+TY1MYiEfpvbBRFACAzUx4LfPTfMXLsFXG30
gRTabMWzFmrK+X6MPcgjXPuBGLJ8bLeBCJybZ3hW3mNM5ltrvi6BBm3im6f0HHyB9dur3Q4GIJnU
D83ABd15LlajpJL8bNpHAvMosLVUipyKcv+0w19R6HgSnzUxpTf1C+6fvQXEZ7UkJxn62hVtRmnQ
zy8hRdrMdZnYxg/iN7TdtjeBpAhUMxkuxy00RqWjIXTaqQPAVvmJcvTDNxwkyFDMXSrBLRWM4qDp
RiHGKEaOh/Vv9jB4GESh618mfR9RiWaoiDUkZNOabNS01XYxuUBDmENnYg+eiQV07KIj+04FQ82J
yjx+Q396/BdgE5AT+UPrTq/uS8ZRST+C1JHXm4zrQeFYMN7JPsP8n/49d1iweZyrBnRGz8xDbWnN
ahZ342yOBhBavRFrsIXKnOg4xYqYyPl1OSFWD+wUNHhjG76l5s1+2jgoZZPp8Dlg4qhnEO9CfgJm
dJ9SIekZgiEGQbyfr8VYJprvpj6Px4vmzA30uVnc7yMNiayGsYFwELA/nC9bVUo2EWXZrt5avhn8
rK/Bi1psog6Lh4PMdQKFaIMBRnv50MOY0WiZviBpZrwQQywUap6bglmHqiv79kdCeYuQwcv58+91
0UY6+0j+3nEU0qYH2OX0xLccyJROMu/SOXmm3Z2+HvPNm0q/KOmhbZinAkUn7z6RX9RxIh2ShuXw
TXEl+Cyk71BKWn9FPsPELG4xaLl5sQ1pdtyrnpOHM+gcEDwicf3JtOrHJyvorrfH5qsUAgPnXxon
C8IRFmBnUAV82ot9SRLCDv75Zg9MtYzRSF16nntzGsN8Xsg+6b0pNIgl7mUJqCIdc5R9P4bB8FTR
3y74+pBnKSpcPnp+beaFxssN+QXWm9IDK6oEQJ2jMD8/fD8eBfdlIFMbGLbcU8rfw3tBmo399O/D
5ITClwQiZpvpDiyqtYCoPGenT0FJDaKY+QfUJpuvs+UpIHz6B2i6LmpAmih8Y2j3wgY4k7ov04f9
uNjINcp93MdKCCOiHzJauz1Ewl835jixA4iWePtQX3ke1Ef23N2C4Y7ogjzP27uVBDv2Uez0d2pL
58IRKgUq+HYoC9AQTUrhQ5jrZuEwPOl188lQX2YSO1IdxUvWV0p+qTKObRT8PjwRwNh7r3vFRTGB
3Hxux/8gAgCvYjHo7bPtwUcesabqFWwoaPzMuwX7MS0d6FEEATYAt5YyZNVsvuf9podkBiMw8FDg
EOZAVh3orH9/ZlJ3f1TKGXBDXKiybI8xAtgzzN7EMCCCNY9GqwmHxYXWzkNgDFGs7IxNX2EP6eUu
newcJopmi1jpEp2HWL6b+P3sGsgQLxc8/35+DbaV4Z4dyFYxWPA33aZPjn3VACar4p+5b4B3EwLU
JtBBXDSiJRtYT32VhDSp9QOnImURsGT9mwchCUGL423Ygv7P2zB29ZkkLkdV62BmZD3u9lwybRui
VrxLIS3i1KiDF87kPZ0MQdRZrxMem4gK6g0xyIZR/67yPIYVCRSVu2b1UvPdJuTLIa/vSt/tbVOX
Va197cJHVJu3gHtjQWRmMBqn70LxgeSAkDi42Lk/VItklVvdPVpTE4pLhH9g+3DuXgGRcU5UNK5j
IntcmJc3x2pqT8sDw4N1Z57MfGb6kHhQosKWbwti/3JNBocEUUGTHp7OMYt3vDuVjgQPgjYJs76Z
7bVK6zwoJKJMCuNEf+dmJHjw5btcV/YTqXMuzVdnIUoY/r8VO7qCUHGAFYWA2Ye2vpOzIgcj/09h
OIbnOoP+j/MByXiv+8abPlKTnB1YjIf5vt6tRmSLSm7Ycb74PZ2A+WOmMqrGaV/eYAgB9nwP5gUN
9q9DoSjxFA2Frm6oqKDPqheQcPy66e8oxw/xGuDB+BZ0HZeHX5DWYvJkSM+WhJp9rwhdfZ7mSwwv
vjwzf57+tYiLzEINQ2AZvEtU2VVXPoWAAP0LlA25906u60mU4mZ45rYTPUU6+HOZ4B3EKCvQed7O
qvoeHJ1QdmvPK1uQLHP/aJQ8ztEbO1PAlnx7gELzJ07yGFNNl7g2DnBGa5lLEUheENgMcdWOTybL
Ozagwgq14c8sUyCixGYVD88vR0czqb69o1bEPIFJP3yj54xDmjntcMGnVmqE5+MR8FDnZo22T1Ol
1kcjE9F5aCg+zi6ri3Pq1uIsCFpxlwE+6i10a3M7A9Z/x+uZBnK6AwHb0g0Tfwb5aRUCnDr46rRs
NM1I8erE+MLI+3YM+xjTuYoa352pY5FxjBOYZp48ODj6z3GwAn8src/FBoLPV3L95IlTGTqbHOL6
kySXB6ZZDsTMmjV6QUjDpFtbuBakvTB3+uBJZ9jTnUqpqrhD0IDuAyq9CaQRXQdRHiVsTQyRTQP3
9aSu2oRG6WRDjgMS9a2XTC8bs88ZajW+4/VY0zXlFtSBoF/J05rdKsBdjKx8IFPnQ6bG+nUV9n1C
/m0/ITF2zV69dbxjqfjFcb5pZ9qneAuGuRaf0/yUKyKN3p1YX4YrGRm7ct/INuDR80tLu183KZjx
pv/rGo4/qEOkSVInnf5Q6LMRsY8WbBgchM0TazxW3l9v0SJyIQZYXIjqy+7Gn/Uv0wrHg63bigi6
2yO2KfxLMAmJKvi0FdvksLeKIuOmN0DKeM5fslfwwjf4D1LyBJwvQMNCJ7GJ0ZV4syhNtYMLuYrS
XsyFFy4HL1t7QEjV81p7mRMjGU4xlX+8ihzIQQczHd7jdDt8wOPv4PtGaEnteFg516j3VTBGqRFZ
E/FT9+YN+W3XGDEuw0i8UnCXq8amSd+v8U9WKbup/VeUEirVdOTblL8zhcb5GgtZv8n4U0Uu02jc
C8cqYJYFsL2xhp/s5htANJ8wrwleE4XLLbWllHg/TlI4XlF4zki36JJPBThYqfBF97rtpbRdcAig
cBo5dl7EBRlfnX1mrB8uPGr2GeBZh57VX7EB6e7nncXqTlkp07w2j0fa7A1qOsd5QWD0+Au4xgKk
O9+2I3waXlZ9e1WBDPMgzLNNhbEZu+PnSFrpPWx+ZtZvoGVhG7yidBQ4qT8qhjrzuxL+i5xnUxf4
ODUlwFC2U9zspFpDcXoL1MKEkUjMH9l52Bd7gQaxDDkTqtwBXZOAF3uhoJMxYpQyobLD77np+3If
NlCgh0t9G9dw67lJwdtb/tqIMeVLi0MCxvyfR5XUezIMIZsrAn8hLtykZuZPwHdqFLp4Ns3e0Kaz
d+0i4hS4WvbJgkR48P0RJAGU8tZ/P1ovmMbAVxs3k/bEYHZ/PKyGVbyXJd2JXpGbuj4AgvwRDbbJ
+C7bqmFRhJtD4SbrwwzdA8//ElLbGwcdi1fGZ8XbHhvUOAARLUcR1ZOExCmyBV+QNs6KZdIP3KcZ
ntnf/WDqPYcEXk+4U3H+cHBBSuC8SErMjSZ5F2AeK7xrYdfNsfPaNRZyf2kJOX0MQ58JG0g4mG8m
15yhEmkWVNLf1oOXrN0+I/4LWrwatHsIuSTb6YrqiLpMqEfOm4Kq73ziaRobtjBtWZ5ExY3LaBRJ
BrpM3HF00D73qla30hzA+dwERCt5wqpsQs22XHTkdzdyEQmZNAvMe09gY0Dx0Xh/+zhfmaeLTfM5
4PnFztWJG7Kzd+dqHcCudC/FQ0UJrqiKv3A2gXdiI1n7x2heyS9J8v55xUI2UO4Gy2kJJQbqSKZg
pJElc87HrtK/Sw2h2ufQJimhfNJoUV0ZHj1buLMxI/blcRVAGGS2teL4Jr7nuCwcPAQH5FvlOMrG
s1/Mud8YL0qWS5ePb/c/u0fUrbq1sjKqMeFKuXY/frp0BtNcKpPBt74EzidO2B6bsA89wbx0lQwl
eCzsDP5tOVkUJddVRZOYyYGf3s3ze055sAne/xLO03pQzLfgx/ZK0Fy1oFzyEP/YU/+KkAoAkVbB
GJ0xfrhRv7GG1Czhe+CejfZ1e9docDHyzckqB+p1yldDx30sHeWgxWnvpqoFCzUoo3VP2183A2GJ
jQT/Jvp+GDM/ZPHTRQl16GtM/J/wI927CWdgFEOe21UwqXMXKML838803OdZsuDKQ0p1B+qWmZuW
1qpDmE5rHSV4k+5SyQp4+6M+veadp303HiE510C/C8ANT2BZOoq0XQN+UKyV1N2Fbry01alRRl2I
tcQZDdK+GbsXdquyzynr8spimac/58j2KsE2HgFeJA6Kk9S49V6W4oIzjWvz3iwy7MstXWQ3gv1l
WXOLoMFLEXqujuu13FNoh3FGAzUUo/KYZ3nI8RkfKINWsoDhXUNxFxZaOMVgoODMCD+3u98UntWt
2YR0he5RKFsavuX6oY3eMdKj7559kpLvtdfEdxyT/OMjI9avtCBUEQ1bIZRBup6EPu/yKQULo5r5
i3W4NH+6AzpVNPdkp9CSF98L3hPCHvMy8YWeihGhiV4XlIMaxE6aA2s5QvEPxM6iHD+4rUM1iEWL
JHhvZzTbxnO8EKHjW3P342mU6t8tN8xtw/7WW8QA2RD1DZ6QL2CcYjRUfaNbOjfILdKzFSDnNbnL
w4MIHxg2anNozyyHHO1iPgsZiyQaeEFTIf5yRlfOHMV7hFh6UcPsH+edqmqL/r9TjMuwxqZAjR9T
Roj3Hc0oJlDuGyECj9HqxN5iS3eUeMcrWwOGTQZcGgvs+3ZeqABRI67kNqpqkOjVSxtK1AkobhE5
YuQcPIEDuaN2A3np3e2j6BQMmzecisWam7sO4LzpEWAO6Hz3Ehnw9y+w3sR0MaUwkjfGXIS9VahW
cZrPYF1bbwzEMrqdsizMAmUFnuCv4UCEed2VUBApSy30dlxkkUrjaybXdOWwHIejUwA8qHCM7wHJ
o3eOjV1fpd4BTbU3KC30DW1wG8lTfP8ke3GcbuzC2eYiRChNmpJJMcem4eQ+4qqnD5Dbckur3hEZ
jDbsfKpeya9xapYMuCCVrPVXME7b3ipGDH6+2/Zj0cjofjJI9NkZOaq2gx2pGKvuJUFjjzBiyWg/
bA2laplDrz7wOCcClkmwdnOstjjlxggVQS8rN9eZ2y0yWVypl4+2JUdFIAApmRRQNjJwO0fxDqh5
nfXS/9Pwdhfy4Q7Ig2ajBL3bPSF1fdD9du9HZxpD/XOfXfsOgHjwgyLhXPasOWzOHZW281ZHaWFy
cnkT+dc9lkEN0S8qOqX6oE0k3RASEzmN2CVeNlvqBrs26LeafRiq6V8g+yxODv+ZQQtPKVKGil0Z
8HgkH7dKmjneBDzMnZ64kZ14vEO/uwDTW1FIQhD94d6lP7GC0Sy+RyLeD3P1+yfGmeBYq4odmvtS
1R6J5nQ2/rBgaoeHbhzO+aSZLRMuHewebCNxkIv/erqf7vuwWGEwW+WCLQLiqcU6PK7KnzgtaUER
PpRtVNGoYL8TgKn1wF3CfmB82LWOhdIIM1itN5E3QiOEkt14T0Z8PfY6Ban5vEU4uHvjQwQIVhfi
KUT1400dl1ITssOaibWqljiUevMw+qVM4tvj7Wauti2tdYQQW2cjFOaDeaObpsggb9Ga4on2wdS0
SlTFOLcmQHygBP9kd8/GdZ5rxuxzNHVeL+KtgLIRRfGq0YfguPdxMDoOGL2e25KgRzulaSx5IfAp
QI1GhbGlEiatGRkS3amijiZHL0lyur+He3yTXWiZNgTGlVO9B5xEAPhEW0C4FushR/5LEDzVgUAR
we6XStDoSl0+fv9/HyEYwxZg6kLAQDpJ2htgTjmbp3bT4s8CX+EThIv3wlsmoLJOD7od6umv65fr
iRRn1BKKwSkidIVei/ColK389tporzj0U1Y3KFe2dAsqXLw2DEe4PBEd3mwVJvJ0jqAsvLqdDljY
eexB+Eo1wUs3rdoQmZ8FFyqijq96FeafFrdd8/IhuxPdiW1d3K4AHTwnwyRpxvzlNJvMtMlLVlw3
7vSKrpmLWBXrbZG8rLkxKF54ibntRb+BURkDcCDua5ZpUiv+czlZdOl8hKuegq91ZimYsdALv5id
k08NzSoxFxVqtAp0VzXeTDTuGuJi2Dtn5LmMppfVIb8WVlzhZ8hCZjR4iuUMDjhGXNV7gC8owWJq
bDkcFfSzUcUoQlnSOY+rZ+pcCnbPGSVSPdkMno8y8AjWGCN89DZptAoBa1QolU1cNd5wOL0vqNlT
F2lcAK8rM+2FrA8AoCWxgwU5O/DXGSEmBzFP1KWGgEq9rWlzx+znfBuL8GHTaJdfJk9ombMqU53J
g4MjJyxiBxKz8MLOhAakLzU1zjdEfJOK2UG8H8VpvKx9AkmMW4c4m7B8SJtVvCrGyDdL/t/1pPZi
kd2lDD98X/h7virG9bmxh8XQ70OMh8nYpnxiJkPdGphhhrtMTyWOVDdVmnapJUwsUjCeBXEE1ua1
vJlXbRNqqV4yCHb2f/lyTgLaAjVfNo3oCvW3Q55vTyM2coPDZawCDIu1Zq4EbkSk90OPVpVOsCm2
+ExSpf40Pp2dYKvp0v4tX8Qd1MjRqgnn9ccVip9tW/2eeyTQBAuUokLrNeweZvGMu2iJjt0g2TXM
owtuzMJwaBnHaQWtMPds1M7BOvEca3Pi1pa3vZObdkqmYXp8zSR9lgPsA3+vnimyy36LkBf934j5
l8MvOtck3T2AePMskLV8st2aZh1wCAxROCtr8S5/wGMyfEVv9M4McD8ULRpzxEEZq7rJMDYGzfdj
WX3yTnehMiJmasgQLH+jZIY0qJwUeyPO7IhW68+j8815HzvRst1/J/SpXUlDVRjSwh7zBnY5jo+F
j2zyUJinGxh+C7ii+B9Vv/n5tCdGoZs77mChuZHuQBwn4fk124eGjcipWaPQ+HKOMFyOP41fEtG5
Zz5mrl2Al6ESoYRtgfKYircfwicoPMaXsuwot0M+4rLddb87FSo5nJ70N8eXA9KXH+nMgG5zsOQc
P//QTvoDVp6qP7ZJ17gLiKSRJB/mnXneiMnls+BBJy9U8NCyKbfOWOyV3OOeVpOTWxurZkltoPCh
YhD12rLZGfebzbrQqtNYKbMA0E0BkPwRewy9Q2UhMAI2wo1SlxAj6i1bO6R45gL4k8Q2jrEvtOWH
kQUD/lyw03usK4+496L+qmSkJOrBsBCxE2m3lRqizFcMtzUDLTlP0ZWBWu0JvZr1LpWZlk2jibmN
Ae3B4HDlbAKY2gT43A1zC7iGW4mrPGvOOS7kBw6YYS4yEdzHMCjX29KFxklXLQdPAoLJMx5oEXlU
fsBeCiqRHQg2K/6AdEt/8qG4CeVStXo8kd3GJKfm7g+m/A4T0NJ7fkyj3p01aFe4jf/JbFW4d1YU
/DN26mxY1+31GBIyEt2bZYqgfigY/5mQz58nEPZJJo1yhAuce7UwaHKDWgqUtunhYb8l2+TrJQwm
yl9Q7NytSAJGvpscfByx+7vdTRUFgC3iIMpcSVsvCVcLpm9wc1oU7UySC6u/mAzT+mXZb/UN0L1m
aJbhpS0dXrGh8k31KBn+mjWOdlcpNemAy8m0LOyhAmO3zchNcDQA72MAWClC4/Ue13OeuHOll1zJ
1xIyqr90UvEcwNNnNn8nl5ov8CXkLjK3UXs95HKeRJ5rc6ut90stthygc1TaPcSfYYIe+TXlrnNM
NMNNaa+C1QhPEWfBv5B0GsCpnl3vHuMITCjYckc7fumXwcWFgY3nfJ9VaAu1TJ/CBrDt5URMMw8V
IyxAoKjhfm83SB5onZbJfZcxt58Si6DLAavg23oIGLk6C8/kvwW4JJh5AA+/pq6D37O4t0t9gb/2
q4ZzBLrPNNKqD/lLWZjcgbN59lrZBt3Vy4x/JMXkk9JXCUBuFDE1UiZXNcYhXkQifyIo/bKutGPI
+IOr9l3C7nA0LWFnxiqCToKGAlJ8cFs/q1895WPKHivWydcQBQtfIhctfrUybOvrc4iMMySaDsZk
7+kvMuMF3oRCzlErDNNxKbqnNpr3b3LtLs/iqqFo68GcmJWTxDM5Pvd/n8ZqsXtaCzYP8GUmEy/z
uBj5gO89HqXP9r+BHvjrGJIpGqxT21AYwlPhbHbiWSfiMXP6yBwWoluDm7/UOVYVZ/NNml6XNzZQ
rG0CQ8aZFKUvP2aOkdYaRwnB0lg7O6RF3r260PgW2ECwqig7i0oWVTMc2FmCSdUnaxiynIILcrOK
S1SnBrYZjjLCF27xLAcsG1GSrCVASq24c5KjiWj8EnJnX6IwlgTVdsV8mreJYo/8x3g46+c3+6Ae
3a/pnSmiiOwKjgBudJMESUlRBVM9QVclVJtWuTiMVAO9Rxu/zlRgbAsElvHUVITdNNe/ieK/dBFE
UJm18RIdpwIqhUQ3EpE1/6RPMN7JzeCbgvydIZx6j5nC/G1zLWdkqM/CE+Cc9calSHH9y13M15Kt
dGQusk8bI3ra8WQEs8HUmq8omCfrwI6YoW8mF4q1NJ2m+P0U0Ndw2EHMhEMVdsDEhP0WRmqmN9Gb
1aQU8IFuPJ8TNkAEfsncjGhSW5HWj3njl7elQ3SYzLXSbMKsa4ebB4X2gwmR6A5SltFP1dbPD9mx
1ErO47m6uCglhpyirafZsdipfFM8RMLk6UwPU1psozftLdLWTulvgRfOa56o+gDV6OJQV6y+78tO
65rLc2jr5o2VXYXQcGB+XUpWwTv1Hh0VnPITfy6IdJWu8nISjNcTUwXDoiB2aG9YnJb/yqaDkoHs
dosBGTCGvLFINTCAmojplp0wWmOksB+qsUAMGcBaVOxBZ5vgT5dU9bUfWm5kuKf/GfBr7SU0Oknh
nv/ZxZbyeuurLML3I6nzyYnXz89kdio45atBT5O4AbpNRAnYz0djALMGBBrWD7nKyUIiHzJ/jwX3
nFb1emy417llbf6rRnK5XV5oXFaKG01XTxC6z2qOHJy2KMPrx/dT+ep0FiNLBfWt0SkkXvpFDc1D
GbJ7vTjXtziJaFe98gBNzvqW2HRzWvWgAQC5Ecw8tVNt4pvgXptPI/klQchh449Yg1V3Aotthw6e
aSV2b/GG5UWv+MRIEB2USNyJeI8ZSPEs/Dsm4yaDuob6jZAH8W86MkSNoRmuAyLL2ddqW02FhcSq
Gqab0EHTlTyRY7bwaawcWs6n+Qe+R+9mIQjUHDReBY+njoaMr9dV4r7lKcWVE1ciWryXZkoc05OD
2uT4wGe/i5yIlL3FvvegBH92G3MrBTIT76SN7yTvO/KQ1i2ciOHoe5IxJkyM7DJgweF7UNr376ER
mrAB/wJJxxTHsORG91uIzW87CfTe6qPI7/KY56hbP7cPdUixZiPjqon1OJodzrWad82fWrmJaMKb
5/rH58Z73iRN78i1g3G74BnAEkRU3tbCwNM+NspdUMof5XX3X80MvSeSTuwzpNECATd37zBX+eN2
iUKbNS3ygK80oQ1ytU7kqgY1ajeuehqbJHhgjx1J9TOjawnmcVTe15979aP7fW6YIsZyVskMiaAd
+bp536+WHWHwSIWmoxFeVVj5bNcSYec9w0WjDvYFfk7QCxVcKvi43ngWpxRwy7EJLH2Yo0AkloK0
5p185eFBJAK/fHKIM3sQ/RM2AlTcN/uKUhINlAErRir1z15X07uyAPWvOdG5MK537owGuo8PIW04
xLUdZ8IUwGTb75KLgT9iPxPBobbvJC0XRCIEvOU8f8uOONRY+holMtwQVLDU7kifeUbiEQd00aXP
vPV2T3IGiUrz7Fnq2Y07MWFm00sA+cLnZmTd8yumzHsvDRTO+YXBlQLZvOvAvR2LKJUgknxCzG6y
a6BO5iCMPIyMsEfTCbXtGLe4sWezjlu3NrNwHoDnq8K82x19T3ckzM6rwCIxF50SXzw0vVHm9fY7
JJ2S0UVfeIsrNbMa2uUJL38pb2yRpGyFL0NIRLIhhUeNwMDaTRYiTwqx5vL96sXlaZjsOH6pcIyn
b2qKjJlj/pvtp6MTVUoOlgOKcfeKUSX7PGqhqVpzTnFofVqMLcl30oz4WtPjq+DR426LD/j1wNvf
vXUvl4JhO1XMHKnFAvfj7fUcSpdigjnoFcQrrIIDsNkcjY8gdlt5g3gC3BhbL7lIQaVfLE1IL7de
nnn6+YVMHw65fpaM2KJ0XtvrsoeSE0EYstBhwAzLHUZICoXz+hyG5AeN0oXLlsufjy3zr2h+eq4y
f7QcldakpOfWHlAE0yP5cAQtz5a3YyN/SZ/ApBmzobpmsFnzYMyIyHc+D5fy9VI96vCGFsbwmPYX
1/qrwqMnUYuQtBkkEZYRIOez81fMlnalxcZjYT9uV8sZBvKAN4pGm+f95CZxAFk5PO4f19ISrLak
jIYa6NM/q6OvPQBp9adLHSpIigG/TsDCw1PC9kFpJKPF6Z/StHvXBevl3R46QaCMKrrUeZKuMc5N
6A+OkiSbNZQiB+dJeGtFzX/fqeKofh4l2cncdljJV9maCIzJu3oZecGuySX5e+nyYZ311S4Tag6d
dPR0ITTa+zo1yh5hfX/Z6PlCjoF6qPuBVmNkYjHj3VwbvG+9MfDSLBpvd25SjB8mYXJsgIQNORfW
Zb0PZr08oCAq/BdF4lvXJA6DesYzVgo4L/kcZ9Kr6boPGb3g+i76LI7TWQiSytSiWQGSrw/9zRQO
TIlol1ebSEIkwi5IXvJX+Xy4GaAV7vAre4kWQ1CpTYQdG5A4s33nWwBMBXdfxaBKRdfCexWMEo+r
Dt9cwSAqFgn411Z7LYCTltQWGAghf4WZYPp/qZ9VGCANzxLrM96L+OYLnJuhCvM7bwk479/6XmA+
nZU1N5OXTWM/EARMFrFj8h4Aa5p53VY4VKCqnelrtvd1uPanN/4+huBqx+BsDt+9rMn8gFAK/ghI
irxWPRnCbZLIjzEPaeFgLuerjXJNnpU5GO7VnLV1tidm2pYACdzmPtaLFwZRoDnVfOxh7QNOXaan
EwAkPc27lJ/VtTtKpfD4BZ60dj7CSUx197GPQ6aqhWAmztJRr18z4J+coE+Fam6NMhhZIEUF3s8t
cGt2BzVpf8MYwF2iq4JsrLXPWWmD1nER6FyH/rEyxoYJ6danTnzN6QYv3lzWhQ3+IS7hnwK/22Xr
LRtkp4XgDeDREz4g9Tj83tSQL9tvx0D43Yn2fGP7rWf8cldKUKfdZtXFFNYAPSHbsMcI9jpwIFnZ
hLBmDW10v2U+Z7eytNAffOFnwB2IVLBGjHqKgosA6RTdC2uTkzctM987nruqZ2+/8sATWaB0M6D4
G5swVjGPCJ8+iF52/pHoAG5u7zTjlWZVC+UOgjJlL8sBVKNvAqGb+W/k4NJ+p68YpgtUZ0RTIzSg
plXV4OZcSg+Y4gMz4RvivlVHXF0YZ/MOEuk+iAsCXHIOE2rOVg7JLDTXaIYnZUBVROojbYg2gmlm
m6nv8GsD/BDR7xiiWXW1YlCwf5k+wHRNNk05NybK/jAxJFI9tVfZ4qDN4UyOYu51aHMyQ+qsX7xk
rMJTNGfR28a3e1jIrU0aMYPHq92QeBBGwaHcK020v3I7j2xMDHEIf+fQXoVmYN7yhZvBMiwSQkaN
TxN2pCbiH1IHjomOnI2lc+zYkF74tDLukVdWxjb2lLFRxSUv0+cISSvQDPir5oi20cTFy6pTO6zq
h4HKHRLb8YXhpO4U1GB5/41B8RX1sZ9nOMZYctAkAUxlkrTHTnuP1Vv6rANt6A6edDcIRLjl0wL7
79z70hfrBAaaAMki72zqI70gR5nZaJMW7jzYuMoySoQmI8ALY0caGuD6kxZd9ozo0ipJV3h24xFD
JGwVKX8KUGb1R3tiuOKg1UQoiLn9gOg6c69vyleJv2L82liE8+BjAYxJTooguWjYdZvD4a3jcHB9
4hmKbqSHbAnakTlxsZ95/I6Qv4l2hzBT44hWHv45ZjQzC39e7vdDYcNMYqVYXb+RvPD6YwJxkZWS
K6dUzNDvJsZMvtrPOFbFIvbrWVpnWsg2r/DME6LZXF5wgT6tE7Xd0LKibOqZevNdgj8gpviMLwEn
FaePSLozPkp+9LQdHZLBuZwXXWOEkqMQ2L+vpS26NBI6860eCqCUu5g3m3hEl+0pjYTuNb77uUxS
vsF68Fy+v1h6lOx7aF8XH6HmPv2uXM9qxzztY1uJheLP08dmeEAApbn3UlUDtfjTSi+PUS23rNJu
tPsWFwwSFt4elUI4jzvXVhhtondWQ0JoYa7MLyRk+/bUGqUQm+Dt76KMfY1fEgpl5kFXO02Q32iR
qWTPi9EnIabDPpoD71RcAuERSwNyZZVm/IRxJUbDW9cgYeU7eCnE/jbDYrdFF4gP7POrxUcgqypk
tryXw7paqidkyqBMtCmSQ/Lf96RlxGby+bKI+remtIiO3wPXf3yeI6/8m7Wdzbm1mSsHyCLijCcQ
xCE2m+crnAh5GQzcstiqHOdMLPMzOoi+5xV1ZjTVVzj3y3wHQIIopvsKdNw1KcE+/kts0WpDV6CZ
6TrbWebQPgc4d7CvY/WJo3XwzczHdofOqNzBRwNgmJwNX6L9mzNb3NdH2WQ07Xs9AXM2f2IYVDop
QMSeoWFy4+HpxyFsu/Lcrc9XH37yZOalKKN3A6j8bO/k0Rqh/SAgWvDq6rqSjben1sD2gDKW7vV5
rsQE2E/1fgKV0IWvKemmotgbJOerCqVW4rnqkPntMbQJzcoWj7pDeA8d7BfwAW4Qpq9mbgSjak5G
Z7nHaJF5xO8VvOWEJiNaVZmXT0LA2deXuxDv0UrHiZOVFAeGafNM9lwfKyHBaix+2laJD3CeXjWz
RydJKLsTE0FGw7tfDG5e+ApdikddtX5Aj677/uXPuZlGu2tbURTho/q9eayDwWbnh7HbW41ocCPE
Y5SSl0fVn+4+B/VyH9v9mK6LoSdI4HgGsA+canUMeBbTUql14HmFr48iS+ysuVDZi0h2IU1tSq0W
rZdMMI5e4D/Y8g+GdLKHr3ylp0tBMjRTufYDfCLL2LeDhovVwBgsi6d5Uhp6MOq8XHrQ+lbrk75S
5yYTujX7DB3agE2vnNykyHBtTlw4wLZTIn70A4Zr+6SUswL+s/e4r+SyWm1AgpmEQbk8Sbt+VeL7
R8cdTQ9JjyjHysB1sbMLe3njfy4ZSTO++Wk3u85nJHNV1iFZO8P1JuGo4QwGb3beljqddgD3iPZq
NjCO6CsClDcZAlsP9yQjIzaufhYMnutpMqEhbeX8PomUX4BvU+QZwCZtczkMWRPJqKEGZB/tA83P
zPjBl8oPf13eiEeSG52S7cBCqJecwDioUXrJNZHu5D2Am0aRSoMDKRP92vpvO4UtmZlOJbiNSC0z
oCLHPA0yon1TjxZU9PMH3CCJtrGo+URI47W0HOSOca2ysPWyqkvUtRR3AnIFkaFDCjrHPvNvkcTe
cvSif/NfCKADkwErEMW8RlH5yuN6RqjkevTS57KqyOUeqUyJji9luMUEcu/UqIid3aJstrp9d8D8
PeOjXHepPn3QPQSfs7icX1236HiY7n+ReZAaJ5lTkjGMr3tspEFUdQYpoZyRC3EFt4MxBZGisVLy
A5bShmNKEKWFiE2yTT9876drI1D4Dji5JJlFCZGmVwgU0n2pSRL+U8e0+YjsFJHnQgEWzQyBVqiy
2fnG4jDSr6eR3sraHoNYbOIS3NgrzZJEIMQieXvChnn1EYqma2MFzHPBguC9z4ZpVEtUFfiY/8MF
K7Bl0iCjp1LvF5LhJDIqL6NT3BYsaCYCPf0hwpQVKQ5Cbqe+V77my2r+lSBeR7WGYiCsJdJZidyG
rKpQ/KJmV1b46NeQiykK444/3G3+7SmshqHuZJClPJw4C6icE9yudFh9zhw10uvyUujli5e/TXIZ
Q2seOleNrYHOs3rquVszVi0V/OtEYRxzydO1WOeXeEFeqpkscfzzTt79Nc226RNcI4VubB2m46oq
mSzc6CzZ+IRpF5ib4kqNBvIjJHbiqOWYNevi/JwwXgqKSTIoZ/7QUiCW5euPnOj++ABmqZvp2gfd
08d1fBPBSzMIC5dPfpx+AQOLiI4zAw+AmI3kLS3SZF9fVyGtmEOOm1CBJ6dA1kLuhc4h22Bqjazi
qi4PtloanUhQswC2qE6KuddJxbMQ9n+Q8PW1EZ4mmmZBUtEEz5YwsKPl1UWxGQZ4WI4ad6bsdOIj
pwCqNxwYvTBbB0LiGbrg/DUlDpx0T8jxZ/abBrFH0bXgtwz7521evGgHuSLHfucYr6wkPNnCIHzd
sIDZDz0HRU5KXmyD4w30oyHTgniz6eTkZXz06MX4498c+vyUAdkIo35eVz3P1peAoGO0cN68kSdV
EoZzYCo005RitwXnePtXUuJorfRnKVxcO0f5DrN4fy0PRb8inE9HJLEcAqR1Z8TbxYIpbawwg3vr
wwPVfOctHlt0xIt/GgFF07ZSZewFhjlvbcplZc1LchtPQRg+dpiXa509LEGoQDBOpDdXR/HNOeii
0xleziEJrADI7ijXVqdZPk3XnIoex3RsOBw4KFy//ChIS019+KGvXj7ivRgUlgXCI5236Jjs/3bY
7ltOeVLBYQ2XihGKh5H0AuZ5l+B0e/yKZQgHe13prfn9QmbL6W0nDm/xBaKW/gVw5thhBSWwC6FW
rG97oDqwwQQdNAbLrPbLAMD+ex+ZDMHRSssNwMMdT1oYouAntVmrOWZww/7175DIJ0RsZx/zSSu+
rUdAolBLV5zqL2vbMmDBXtMg+26VnlNsx3t9XaTZgWKjhi5+myyMSnWs7MOj4CR3Ev5b3I/DLJ0p
swTIidBcFwBoFKkXI/LvJjYDLqvlCeISQH/x7MCbrPov1Z+9yhepXFg63r7LBODaVAKRYix1JOv5
oNKmoJ0HXalPp2/FFF4Ahr6x6G6ViAEcoHdAIaqNTWZMUkFr3jAegMxZZnV2rbTOhyj5E//oS7Mj
AGUkOYx8Ck9WxeatMU1d++xlQsZ3+pnC9GTzjNlYM4fmHNWJOFl4o2K7GStoUqF02qOexBw38teo
UxgyV19/6h/ji8zzSPM05NdtPtWKkVT/MNp8xOvlHfC2km2sRK+k/LsXxUBWrx0usZ67rJMjj8bG
Dju27GkBNQblJVWzIvCPtf6tgbIZXXPrQ1kv1Is3M/kCTBzjRuwTovVjKAxiXlBGGhGMXCf5SYfK
R0siIvdskTFSlujRhP2CfsWQw8iYsEvqKpZv2+cMMOnO+ylHxTMpKHKHZbXW1ZP4z1Df/7Pnf9Xz
PNsMj8qXb3sx/F6J9XwZHuM/JwgwkYQBzifUQFqrCBqWil/wds1g9GVsCmmiv5pJw7L1K+w+fQFg
+KE8sJ5nCq68NzkRFiHe2Eg3PNEQGzs5K6fyZXP+Q6cpZw0EV9OI9syBWwyTCe4sOzI7c4WXpqMs
MvzZiFD+uvtK49I+w18/pGwLw2wCHqIhXLAqTXCYFRch6uYKgBb7SFawl2KcnNGWeNw3yc2YIwKK
Dn6TpzC07e2vseS+CtToyu+uxpBUVa2et2v0Ge/lMD62qAaliGbLfQ4TinBwjbere37e8Aens/Ww
LjE38WKU7TML/zF1y0a+opo8S0E2yHy0ivPkf/4tSOTvkqOWw+7YBooKzDHpF0LpMG1xonquBLpF
40TLqmZHwjeMXHuFBeCRFY398jOx4jreRPIXcs+FDK/HT6KwK9uPRaywX7aGUpMMqhWP0tU8RkPR
Bupe+3Y8UV5/IPpGlzuTE8WCGJXWWEFZqEyfbHhBXetIBiLGS1FULPL1U5ei4qum5pR3joGRBYtt
41qKBZdLj46CD/3dFMaGynxmyY0CM5cvd30isCNkuZGelBzRZv+aooNn2Vi5Sdv/Rssked4bNj6r
OGbRXtEj/AUMtVCEdpaW5uDITnWIZaH0rLgRaAPHw8QuvKiX4dA5MURVlH1IYoxm3xM1w4t/SWyh
+bXkqeQYRUABvg5XKKO6bruOWQG8OQtCEXStdSImkdnQCN3db1OJBat+KEPoBHBOM4f0kRzDEgs4
Ap/8+JjvTqtLRHoX0zWcwTYZNy8Or8QnvSzl+X2HBNA5qW3HbpUdIqNuZhU7rveiQVcq9Blcs26M
llFg3LhlRHnQYteato8UYtuRIwlFVJ4TnEXC4oZXYFgUaPh3omSopK1nKsFl22TJDFKtJy9+TJrq
p/Rfjj8FD5ZgZeo+7QoK7mic6gXnBJMd0MlupIWriZbOC5gVGSckrmzH4s6+Rd9ToiCy+f8k+WxC
u9AKVu7kqBXdoQ9myzLcxbqBzx6mUoQqUj7dAsLJnbAYyM9VJ2R0udcPILFdTkRk2L36nkeRiodI
2b277KApkmPC/43beQLRg3pdQcPcxZgyVVKPgYF52Pnste+E33h23jRVtjvlLaX6ckWeDhJRdPXU
58jJN71rQfATyj1RRT8kdTA0OwpjzF9V38tExQVrlO9hy5Nkis5MJPGke6UqssEx6EwauyNHPG8e
dLhWKhUS7O2uBHnLUwLJ/KfyD39plId5y7kVrnXWfVmOyJdwpi/nqRrHI9az3+p7UWbaDQY9KT7x
7tkZnZbcV1k4o2g4ggX/AqxSI3fwZvtqrQMz7fBZWigSj8ZzvxIQNtVxeozRG0Nptcmj8T2u0j8H
bMpUOz2tqCvGrw6dyb1cwHHh0MsABnY3J0a5DhAuVeBJlKew3a61i/L5vDwJvYy+QSqLgB9a2yiw
oClfZ4Z1dDEtIwV5aGPSOhU/+eaXI2k7zkM2rAStHSxNpXFKeKvfA/S+9hrVrXbp+RpuKi2dCj/X
fEitlLFpTNAc0YO30A78ZRvd3AWlvuXvdF33O6rIax6Sq/fTny/FB+YYQYhGyllYDiLssq3BUMI7
A2SFXdpz9JktNKPPcuCqAwsxmVfHCMSU/nb1kIvQhzRWT0yMfJzCb8xRZ7u7/IHYr0BmOUKZM0Dy
EjUlGWDwQGb1agB/ENCuiChkbLfVRxRURwHPYkd89iSBa5ZQ89RJlS1pisydE9oxoIRtYD2yhR7l
ImlgzBXsLPr5VoFQzacLEn0OWCYqAbPWkRgqO31tUL7r5sc+X4VEOjWnTZVO/R2PQ1ZVVlF7PBIq
5/FRCiW8zJ39y9sCZKTjpdyxfR2S2NwzohwxYMvLgxzQxCd70hU8dqis/T/Hem7QlDlMhDyxhhQE
qhErpMLm9l3fFXNJ4KpXxCiowcW0iP76qHnGKJ6yI3APhGCFG8vwZn88BvcJoSNu4zM73+Djr8TO
O+EimOP2j34QOq12TXAwI/UaiAA6F7lAD/d7ZsoFUgAX5oX7AaMQ0arpcqqaF/HkBrTt6M3xnHh7
hZXueeBr+WkcWAffZQGu8eVuRYT9Ffn+ayWM52y4Qv+bX3r0Ng/bjhqi9NNcld4ANWiouzmzDtGm
SOOEHLOn7QE0OSMf4aZcs9NE4CaTGcSmysL86kk6M/I2pEHvpAuM1Tk+N+wTY39NZx005YmWfrLL
JOj2vhyeWNLz9X9lK5uENqEZSpHbnvbQuLxLj//2czRTi/34XN1I/aAuDdaMffJZQvtNFbHmeoG8
Ytx4ds8g9L1ZC5MCQxXT3IfJGbcPMBQjSXU/TF0s2Y0uFhTnbphzZZ/El3qBG7dZXOkL8pPhM4LM
GKTVbZrdGZg7gIuDCy949MuuBTQDd5JzzhVhZ4v9INksROm5Jf3A1raV2Hj4RKepYn+Woq1yZXf6
OjS83z6PlNMLn5RbViJrRaXcHNzn/aFsY98PGVVc976aSrgJZTm02UtiSBEfh494Ot4TNBefnOaO
DU/4SUzpQpumzDiEuVdjJ/KUhiz9IXj42QrBJTKPoBEYgPAr5RLl22pRQvD/aSo4QFDwAV7gvVpN
sAaZmPLltCxlwQUOTYarV1h4KBi8GUyDmTs0W+FuNoi65ih+K0pQOq20zGVT6nPwo/SP3yJcy3vX
towMkuHa2Mv5LFgFn6W9HR9z1/Uqf56y0XIdChU7f/plGnqLj9jcNYIhN4TcFYWHTQAEZYiOQKvL
nB7QO72Y9WYpgMlWFhEF7mF3MHCRfywbneVSGkcQ6WyS2kmi/808SDCWOvY/SmP44vzgTzSXNreG
C8VNPugYP8BWfovf+x54BycysbdXvKPDhGGvRgbZ2erLvH1HRtLpyJEUejLt7h/Q1Iuqdd5GO1SS
+7/n+E3Uj8o3Y1M1cJ6U/oMNOXsTl5RXTrIjLOUjaGTJbseLfd/FuajPvw0XUVCOI4o6ftQmsVyn
yMUgPlgE3T96j+Iz2jaZf8fYfcU3XBu1BTWZsc3NHBNRczVpng8n0UEyC9uP+6PiHF//CFWzQ8Li
f20tey8PrQJzT6KdpkwVuOye2tw5t/cPTigHUZP1AjIlukIYl/iuFN4bGs26Z69QU6jdjLQgMiaf
QX3dsDOjvMnFrs8savRwd7SetijEh0wPx+R1mXK4yhV3yAMtLdgOPvrmOQeqDryWo7ighpfLq8Yq
NrZzflkd6RWhIZjptuJZofzUqgBxobHH5WmhdxXWBU65w4ETzxBK3/QGrpD3nOLVo8sWAiz/Lah1
jZ4iRsmWv6UTvxqxzi+H/msN+31v/5mPaqBWmLhKwBjwwQ9JqCJ9w8N7Kd1LtvhMYlCYfwx/phlk
lGhcF2ouxQY3i8H7zY6eVrtBVNmLy+x2yEDcThSmfSfMAwgttRgTM+47E6mXEoENAFFqmI2Yb2aU
O2l4tD2ZVfnP6u3W18gym/MNmqFDsWJ2i0gDwW96kq1UYT7RR0RB37Zes1tBuLbVnoTLwSFkfq1O
tS99STc1tQXWtEysPtgvSNjcLWc6IyGDJ+hkNK+l+geIsBGomvKu051uittRRpSpo++4tMjUJPqk
csoXp0N5OgoXTGpfXo6fWbQXxaS5Zqe1kdhyte4U7F+eFSP7PBKUoH0gk/tBsC7X48h9NY7I0kIa
hhKu6ZRtruRjXZCWP54T+sCEZ0Wa9Aw57+WSMNjtCid3gVgsY+gNanxG+7DKGgy7F9KtbIntWjHe
ucSR+VQRShYevwepGs+zs74tH92xVnU6iDdR4ZhsQpFC1w7e1r/a88w4pw9kANN0xRo+QI1YNRfw
hIYvl1kavngBuKi03Aws9EBoO/+/AJFYWATWO3UcmUFmmZzOpu0Rs9TT+WKBoNAYXCCdQomyxBHL
0MwYDisifgPwTNwU7YfWiaVGjZd8c1IdXawPz8GHSGmgWCz2Nou3I9CedBsD3bfZ/bONzJq4zKuq
wUcWXYwqVZq2fma7wtpzA5g7LAVyaxvK4sYra6L6+YtBxx/dyM8UHAaTgsUj4RTyhJBL9R8A9ZCc
PuiFk9OBKsdEU+oUShRLgF2UUB9XsiBbHl63RGnnvVTzXDHA1f9KYEeS7FTb7Bdr/F3ihPyuaDme
8+hzvuU01htKbC982ilQAF2ptZn57Q+gjXvlu/x5m/fGATBB5BXMTbu8jADWB2uzgu9WQFQIEjqm
Vc1rKUwmY9EMOmI2FWOlOxisM9I2lPeTX/GptiRp0otaM5THPqjPLz0kvZU+N3TFPFz/etNsLSGk
Ynuob1yNje9Fjr5RRgsl5RAQCGFg0DEnJ9BS4G3rAzQV6f+t5f+jaAONcjRj+dEjnHO/socg9osh
Y2bfefdlo7DopNOffEwNQogzRqREhjSMvORsDS9kl1N4Gf/uuzR61y8BPHy3ZpD1WwGPEu4ZFhKp
m8rKeBC2U8DYV0/WiR5GRnv7aVf0ZtTsmIXo920tT8VTzCULGEhur+Kv/93c7LInpIQroixp69vo
AVGcythlkeRQXC2AGfAy3s6MOb0+s9/b63IwJSJrDIL888g70su69OM/j8NR7/QWGP+MbDrO/m6F
OCVUrHgE638smWblw0Y0CGzAdWphlBwE3lW8Btn/39DnVpLx5k3AJNej6f0aApdAcDCaqdysqzqj
kMefozArNrtjLnLSb1TN0/52iY6/9kFtspoRBcy1USX9ULTdr76qx0KrKeL9njcjlNV6TOPgqjvC
y7pTksUvAqO2EAa+8VGcBLYtXvJ9kdLBVxqzrp2NV9ydOgA+AERYqxvLMcgQogPaW/AVLByCysfi
EVe/h2uUL9aJi7pxJ/5l5bbHek5g9xZwv8hMG4ZU5yks4CZdLAecM8TEAlQu6PXMPhcoKaJG1vXC
Qwc1dfosAGM/x4DgdLE14cAqSOAwTCu/IpNsiqJdB2JrcNDFsiYlkQvAi8Mry5vFV2LVYalP66AF
/1+6A8/d/dRvO7+kQojd5Yoc6A/6i0ab0nWut+wh2PRuxzhUKC4xC8o72FnsCwpvI/vDcidEhXZ9
z6/Yb0acT/mlvUER6YsfPbGhDoVogRlVYTjHIVAtSZ5GbUgQ8LTFhzFgE8GBz/71HN+cQvYQX+6S
KhZ3Nw3kqIM0i5YMZjGcO/xTnzuKASk2t7pLeqlFy1kbrBBDQKddWPnDM7j6/MgghEHKKrlOgbux
ZcCmgDcg1Us5OGrf3U3FJM8xqO+mzcnJM9Dz66EizXXseNuA9hMzy7aRhyIhOvXggg0rOt9lJwTu
CKjoQvXUTH/TGTA4W0WIMbNLz1B4mrxmyk/Zx0IR06eCaZtQSscSX9lW57j16uQ+TLCn9uxMgUAe
IYdVfXs2NwlPo74Ul94WlUwXvPvoqZl0hOTpyEB3rKB0se4GHGyO+HsZoxp+gy5owH72kJT7xd1k
JqSU5uPl/PKt4zkMUakWC5djcBkjJ0gSm+cnklFnzOSmFjelEAmMaSHpwwGKgLTvEE9WYIOJUJxa
1NSOsCirVLnmQD/5aCLyxRLIJ13NxlvlKb58FCw5+ZsJAgIEB0EJh5pTrDD9ai+dkULBtJfGECjR
ptCTLnH7n+PSXTCIxYTLcgQt88XWQRIp9I74OFWS6YO16iJezj2X26tSd+d9Y2xv9C0jNx4Y0ZdD
lbm5tPFubI1buIRgxLoqGhbB1dDTmOY8fOtDVp5/kTNrNRPAkvpMhmXT4ireybliAgRtOfWtO8AI
I2FIZQd6/4RZVw55iBqi7YCxBQfZZ0vGVlWXpFqn2qB3aANmsG6DQdlzXZvNO3QvIulGziTwUPaI
krUJ4J0R2Gmks8tug/a6pCKPo7EA1sX/bAqOuDAwZ05c+H3fRR6cSKT5eu3TbLxVOjRVY+RYzSjp
ONQS/5FjtGJB34CAnw80MIKcIQZYeFyS2rbiUmohB1ShkhlFgxYebojmlSzfqQrb5bdmx63Sc4PP
arIJvpq+xBRStsbAzzDzKjBB8EK7SwFCcQpBQ7lV1AIQAQo2ajNjRlTVrmTH3C92kWuEWvHKudVz
h52Z5853gcGHe+9eqyAl2Ie4y0I3kPtk8PAvgKvb97ry+W7mb71Xtkw5zOUxmg/fks2G2IK53ljw
BvOhZUScUyt0d1tBd8nKUOAlmn8qwH4t+3D0I0hXV7vzpHNtjhYo2ZtmTZycU3wORpFz831yVtZv
MPPTyYrf5b8T8HUmGwpj3Cl+DTKacqnSrBxA4rPii7PJcOgAtIisXJhWkv0c/JP4/kQ4gUXK3r+7
9ROeSi7AFpxPOxtZ+F4Wna9sc4JbtIFFltZOx+Kp28fy5q5vQKXnnnKb5bFg+mQ/0npNqUgxxU8q
3lrFM81OV2mnlaZbMIcmVRvGmpZovuFBdZabI1XaPVUO1QSmolQNQN4pzDVRSGttcHuRVF2nnZTq
KAmWFOP6jdm5I4sql7mKbKsLUKLQbFy49aXXKD9tCIVCNVCD0uc344vtBxzkY8zuCM+3ikyR4Doj
g5RGnd2U/mTZUWZWYUA94rZsDdnuej4iTWT9TGNw1aqmupfbyTYhFpRwqQIq5F+y2XO+4ZzaTOQ1
7vfrHzSkvwRMcIQQd9r1REOBgGBBe/olK3rXIuBOGy75XINo+IRqlyabAIIHXBF8IzPEPPwEC2eo
GjUkmqowBxq+/3YkoUzmLc+vIDS39P4J3s29lAzJ8lmCE7+hd4gzaaW0HrhbLQLJ4j9bLv0ZnexD
cOrIuvVO4L6zCmkx08LS6uoZvMboAQqHXisnUD21bEXl0J2vrik3QLR4I7JULFM7j+x4lyClSQVq
JQqKa8xIs0jMmgHz2R5q3J0PSwI+DIuoWnJ9/cffp+ESg/v/qq6ftttTVf+Wl91eNUtOYgF8ELZg
PwwC+us/3NrA/xNWFI4ZQTJdmasvPsmvOFOIU654NdD/nOZGxZ2mOo+spQ9ESvTPCgWmfKqvgA0f
Fx30OYGi8HzAAhuSertmDrYtOVAYm/xs9lzxWB0tzrBg5yHVitNMPZlQkDLWp44RC00s1LZuPLk+
lWRZ+lVGLrG9WRQ7UgkEMenxH+QRkzYdTrqPU+iSWjDwEwnDIWM3oItNzDeNBnu5x3XSnTHwmqxz
XZOOo8dSB94u4kz0sjNaLtWfHXe4UvxzOBHQ26y5eEnnt3Y5WMIGFm9IVGyAzuDkhlW9YzXxlrNh
Pdkx1A7J6M9ACg0B9EGSC0AFMtOGHuxOCsSgh4QqZlv85uKEEVAtQbX+9tCkj4O/IWj+BeseItLN
Luea2PNnPU7Z8OlNHNRPhXNhtKAoykY6/WOQGo550GpgNQNrWA9H2THIv65CWFkHQcAFU/YKwNuW
j3C4r7LTeaguGGhM9OVUuwMWle7cosKGrFa7NISf2K33ctqvfeCnztU0/uh5W/hoR4+vPM+CTlL/
Wmkbuf0+ARdbbecowYjdw0BAT2M5XeejcPz4TTekUBtp90jBRtRjghu9yITSVSxIResLCG3ADFhc
Islj1UJlb4FrbHl0aDqzOXKZDovhhtZhxq2vTfkqxwK57Wp7YEj9Mt3BCQsdTdrn7rB12keTqxtz
CyKXzH+6JNTDUU7BORLslAbPWnish5n8j/XnA4sJiMy1nzImX9heVqMnLlCB5Nyx0iZqfbwcc1Sy
ahrMGmgztW228EbpySstwV+mWTClIMA6X+6Pi3oVSLKvQ5Wnxrpmah9rrCqel5PEHO7DjgPDdJQi
fpzBs5pU2ie0f+F34CzNxId6iEw6Ev2pSACepHKRag7mZcd6vcBUm8kYNUosUJHXoTM+aOIqY2yC
zcEjY8vTHCJJt7WtW+/FhQ7qi2r9U33I8bDVrNUmsiJUeKYUPaDgWz6ehV2sF2dMlTnZ55OX7om6
uziy01egWBf8up2lmHOMNUUTGyuqhtuekFaFofGdwduRCxBcx03qzKoqLxJOF2FPBX1Eb3M154us
fkOHXZHGbOs5rbWog7QQGjPA+gcRJOl2AXfdSWS9VtBV9tMoq+qZaSNW4aqDaVhri7XXN/kqXaSg
/xBgnJBGklY4RNTNLPIHYi3mQfId+uZdtz7Fkxm86gCnUrlZ2A6fTzUIkXpjO2I13is0PspxwoA8
zOb6s25HlmsHRqmYjOttXksSLBVr/UdgbnyfXaKvulFAEbnchsLwd2WNUgZvbbOLCOGCfYKlf7pN
IXa7ar72iiZ1I9zxEq/bl9ZR8BZDuiyWPYiyGM5cXWEpu+4PSth2GfiToSTZxDTGR139gEGUJHhn
4J0fZrqCBaQhQJ0i8Fxr6u5ppXiJLSIjfnVq/IqR4yaDCUjTAq83fVLB1HoNUWcUaVoqayBK40YT
KzKRlQ6sehnGm2H36WTgZ2ftUTXfaP8S1M0/SIiAtye0V1iNLGBR+7lHMFMyyrbW5k9ZkQFgmsMF
KLuV9dnGPUgHbMahvIhEmFqYQrm8uifit0nOEp/3l4ubfFJI/8vzHZaWN8GQR3ajHhJS+sYaRoCN
set30zEH6z3eHuxIFloSUic6FnMLwueIDTXe1h9C1SGZUswS43PtFUBrYp8BLRYtRO12pv+W8cfm
DuGvOlFZalMlz2U+ETPklYD/EjoXf+hScZ41C81g/YcS3oaiQKt3J/gU2cvMYPCU16aMwVTQ0NXa
vcU+u+/OhF5+WWE8Y8YbEvYllmZySc+JLpOTMrgs3GM05sHcZHzi1PCMu4bBXLqo9+wf5UF1QWkb
6IGLl7i5GGiDXwif4c4HxP+lKWHffOid1eQWDtvuaR2ddh7ID+LZ6GEXe+lOW4KZo2OUzEDr8uq7
8LtLDe0WsIYJXtSn0nSFN1mCXaNGzfAn85B86cdHf8zwCT7x8hCUVAlUgTaBpMBvT/fgAB+g/OHu
G8V3EBDqS59e4IHY0zxkVKSeo91p7lkDROBCrNSpMcnYEw+IojG0Cz/bUd1SVzStIeoBZswniPKr
A8Nit34Ixs01M5/dadHqINuiLjj61ZYL1l4dsL6WvrnwlsdWkm1wXBTpMESt04a/Vo4QAwzVjfAX
Fe317/lPQnIA4wOwHox6JdjqWStLdIYL9wSUSxqkQ0uISAr1pDyCjRLvyVxQUWLSUZmvKJkoxXNh
jPukMTAazohUqfBWM3ZRAld/qGqgGas9VGq8e1pXn7P4fAlOrI0VtE08cHLrJjeUaG3vDIdRRoXk
7v8MwYD+7Oliwo8A3m29AwgkVvOwYLjFpM3/xseNlmYKKVbg56LiSYdhvtgpQaj16bRwg1IfjX+R
k46d2/r9CjKPXqN5ngOIgNBFXVf+euWjZO13wvlB0CWs/SkGKaVITG+A6O9lA2zQbzH6bDZ9zFQx
vJ8KQsb8eQKRJivL6e2yRlJiqhEcJozoNE1m88AKM6qE+Jt3iqsOvLyKpYjE+RH6z8MRtKszx9zg
XvxfXW7g6lEIb3mEJvtSSvc86EsxkZqatcg1eN74bIORtG/74MeDAw/2EFysfUUDwHEMgWIjzRsJ
npi1yr0RBqX5nCXeihtZ7D1F8O7FUquo2g247idTNhyPEE8jLWO5ZaauJHhvwwvJ/O7sFYHo2puP
uOyOzrFzkU3Ly2dCDUazygkFC9XWYo+99/+3cco3KlqB7Ki3suYzCMrZrvFtz2Y/L7nYjDOPqy5w
jVw+hrL7z35XV/+WLz4OqKy2L9CIlJW1i5+gIFR2dM22udNQXT/xgdinTFL9U6SdkGd2v7qTmmzn
u3yVpPiuMw6SKOlRSlTj7wSmcbWqtXqI4g3WnxgCQWaCstpWwCkJRfpa3YiEqTtwX2s2MHndf/Ny
QVVfQEWN7EbnJ1L+zP99LQJzXaqABr+Cgxx96CB6n5fz8wTHf2x4PJ6qocaRjYvXI+DD79fliWv3
54VrxaWBEE35VPEv/fogGfUTHqrtWSVYra++cp2Xipe6DklM3nPPS5pyPKGTWXiBpdDcCGd3kDMB
dgC8BZKIwPYbB9IQRxEdzE2VPS6EYzK6rIIArNS27o6pPkO14qpmCBh/QF8XQ5gm3KCJwrRMrO9z
c6xlFEE+5ds17ZbbIsHloFmL31igOlYNN+7MYQKHZ0Br8aY3LgRNYTBCrJE+yqwZDMNQ6QpMOsvi
C1r7rCE202ZFR715pfHnS20/LWnrrGoSTGkLx7IWDesk9VQbrfoOoKw2x8Oek/KETXkHiRrKNUwl
gyxeHaGaYi1avlm+iPaTOWas3N5DsML+4KOqbtA4VE1OGfO9ZncZDA+JrqHrcwht8yPFkZdFz7df
kndETeS+hhMhY27Hg1sAwUocapklA+EexYiae/ofHVMuCAfqHm48w8r21t/iNriG3iWztwOljQn9
O1AD/r143FmluRfCOK/ysmVSn++lzcDk2UmaDbBVgb8SojsOacJavSUfaMukrvcB+ROdqwWfTJtk
HCwxaHVPGQy65fo5VrgHu/J0YC6//6V7jvXXecod19XfKLASVkRiChb+f1GIZZKmn3Z3wMB+Tg+E
Y99fGx+4Y364ltC7l4Fs0E6FJcueH5KvTAoQ7tnR2KU5QiWJjUwc8Q9455K+ZsfVyIhlfPS9PsTl
d5m0al3Ba0z3lmpuThrfyzHa1DSVfaJbwOxn6dexD87WitKETZiiUvP8U6M+06v7N/KCj8Nxg044
7rjyJNhdxl57De5n1tMmWOFZofCatgPV4nD2pCOEMQ9DIw9RS519bC6tqsqh1AaOi79cFVx1NCAU
ifeshyogZ6t/VSJ5dqTLQKGzFpTokRiW/yS2DFSX8sFRjdTBGrOebdIIh5nqjQ32qTOVA21EHo98
S1QmrEDrT8o7vCd0Hv7NpmPucD/VX+PWm3eK7ffYtnSDc46KPR3DYY5iszZbSjqx2Jx20vhPQzWI
af8f4HO7ZsyXhBG88tt1qCFzdRMsjXw0VjtcCspaLcj4TvlfqmsohdNuo8R0M0sTg8fNzSEIItmD
VC76bRHrbh8txs3759qOO17JL4EoiM9yllk5zvcrAn4tVq2ojJ0rDaDaoa/jw7uBU5QEmiOzVrOY
3nZ0wbyqa+Mwzm33fd68NQ02Zn4DAJQrGKNLOEOY7HgLWFYvFLMSzR6AnbuWcUjjvFSyNk80mvSl
JtEIemLYLX4dFkgsTCVLLylIVF15NCq9/5iBA5500jkVPkpsySg3OCefzXh676AXGlf4YNYOEKdl
1MhM+nR7efmwrcEHS2tCRag2zIF8xelHY6BPgyRimK3QChP8SMzRgCUYJBYKrsZAQU+Al25zgmmK
Om+6oLkW7nnnEgl08j2jB3j0xSjgWkP/yTL656GQHxHvSjglcT7DkoFe7cDOeuBVB4wDrzSNzG0l
PBeZunw6HGy4x336Rp8oqestxgEws9DCEAZGP+EXFpFR7vyese4P+0rilB2h6TeucZeK2woOvyZ4
iB1060FnGHdhoxe+9kZAP26vEnb1sYKTpKw7vWPTWv+UUs7zHCs4nXTUCMtDjJ2nduj15IxS5yfy
jqkA7Aw4rMkv/GiFXML7BdDj0d0JsuwoipLTWNKfakwSyuc/1DlTDnPV7f3UbSQ1co7aWRvQEJdB
0Q5md4bkW13WbgqIQ5e5puB8Rr1mYXTKMiipVv2XEgl+vWnnUsD5RxF6AD8wbkvsGUiZTwm+d9Lx
k4E6tn5JiRdX2fXjikPLELHAMoGyCKz3/9ykXs+Ca5knq1iI4/oenyvK7zLZ8eQ0VBU0dswL519m
C+oO7HmpC2gXieaxiZjX/YGSqFmy4nl3wXcP5//ftkL/KtGPoOf5TGcIDT8zFsbsEiYbeu2fSumO
u9t+X0TzNlFr21nJlVDX5Qjk/aPTC156P3wcX2YUTOdhuWYSONtlo85C70q9XTi1Pr7jXUQlKHpS
Lau1aQ7f8Fab2FN4Zialn1npU6uCyNIndxwBX4NID89D3MOU/SyRZzHNv5FXbF4J/Kza6/CoXEr4
xCsQO+Jpi8zU3yf5uLBOvb61sR5WCAW5G66IAGvMM3IW60KCxdEKv7cAzN9Z0nVKSD4TAjvI1sHk
FmEssYGr6zW32RtB3lqrMFzzy68jsNdgzK7Xyt07rCc3FsPNxyL8mBzoemqxNJTV0bccBhNVEqqb
mgrk4B3Yt8FbtnJCc4RewSrlAWPDa9G7dTIqq8hQudg35Dz0vRhapAB4Ovb3fQHPHRAaF52kInA9
TTBj83dQcrOJeQBanEiTDF4p0CQw0nfg3Msth1sbfc1Kgndufly1/kSpxfGX+IEor+S1wQ3qDUD+
+ztXaN0BZXkHqBeVATKb4d5FolrMvE+wngCy9lWg/4kqhphBBk58sRVkv8zc5kVAN9j7/avBT1/J
/YB1r8t4pb2vguh8J/1uV38nlyK4tnTCP04ncONe/l3COvvX8lDirNylLifFQsuqLT4LEQmsqz5l
AdlSdx5PGY6MgHeZh/UoLDW2PjtQnqWnPYNp5/AIxnbHNoRnrCA7xSyRFkeuFk7jLCoffv4Pt1tw
M0F8LPI4dNEdj4+UtewxYX9pLXf2sBWjMYhFCumnncVb/lhiAcA+Ut43Sk9iwXm13ezFcHGS101j
lB/qZmxeT1xHAQdVMTrNL/P382m5GAwkduxusH9erV9WeYB1B6KlfIRSZAwvoAmsg7HDKnfQDbes
hzlnb0NV3VM2FYh5W1ZA6MbwksTl5vvwPAnAzcEADsnivzMDbHDbB8oDDr0V9x/Nz4l3UeKxH7QF
8LEneAxqEIu8C0qEpjp/vbhI3IF0Y3iQirBNdIWr/woOhylD3kVKsWRn9cEn/WlMHvUMXuBJ7m+L
OKJv6FyJCD/ctXi8Ugj20DL5veC/LRFzYqIjrGN6c9nk6Oh9+7gj6By0BImdOJ1k5xMiTzZ8+Wak
FEg/Dt+JFXPqNabjAgsyc8kFMLncbC9UEU7BgvzSZdKjRrZ27blsmlkMsn+lbN50KzOsY9a973Dv
kfGKCbF6ee5saJ36UwVGQlGss91esY/kzhv1YO1D1gV+1xgEfXna0yd07n/ylHWiSeaM8TtDh6iX
hpV92/ZaOwtD7qMi/O/TYSmVfS1gOmBnedAGuA5boj1MhKVOSAlJAT7dzAqc0O/yOk7YmnSniiZl
cjros4YrPmmGopVKtcdEW1DfRv4V/24ywwM6f6z3XhvgyNZzcAvqmfhtrWMDI5YPbB9FlspE8+Wc
+gZx2PwQ/e0kaB2Z91uwzsaEIJUERbIBuf86pT0k+o6qqo62ZpuGycq6qJi47g8TQ6P1p6E2MlPQ
ykIp63/Gcfcid4SAtyyMI8dOllX9fzheBIte8uVBqgNJfgl2aqK6MD1u506Ta39fKVPjQwk2Df7T
Uex1yIxs9cTUTT0wd9ZA+tVaRTWQicSROsFbUIIWm2gRejO1uJ1Li3D1/ag7Y+9LK/LPYCTwrEzH
IibPOxJ32iFmPxYUPRcYCRslpsr6vWm9IlkMLrYNAGwavgokIL279dCJf5zy7gKqAylF1dp4Nsf4
YUJgGPXT4iJxullzcpD8gsUd9Zc/ZDoe84uiH2Aw1BKwibUNHnkC8fLJDTebMXpt/3vAh8aoYJXd
bfGsTkmHaMUE0SSt5cmOxf04gBE/k0rwLouxS/UwbK+OkTCso02DP752WFpIE8mQiwaJZWNEkeAs
jxuNCDXSj5ZX44IzgWCrgj/butcDnWXp4yfTPtE8V2phh8j5504xm8HeqKUBe4nZeDApMpQr/+xK
Av8h4K1LUfx7ECBue32ICGjEHds8WZmy5YfSGN5wP2CeAlA2Zc9LgznoppwHsewvopBm+ttp0bz5
cQ6B/sugYUKwFgDUPq4dD5SafYQLOWxmkSrKMNfb35MjG99amv3L0zrb82NIivmH5XbzlP+5hgKH
YVieol1082b5vPhA+sgZTtUrARwnvcDDwW9OOwEk3G4fp0wFZyL8Y/yDmQw1/5TcOzYI19iHDvYS
aCjqXLiFi9nTNf6W2jwx8ikxCaHfFVFL72AYVXOLI34pXAd9jOlQbBdOyNzh02Yu9xr6QkY3OCBc
SVrj3yJkOWLfuhF/Ld6nvbNOPRih/6wwNeOdXWVrwaoKfmmwJ3k9Z2Px1UURz4DCIjXf3FHz1nnD
PlrPh0ef7I5oy/CKqYc3OstQLBnRlN3cSfPp5m2IMhBCiMJAz3k99Ki92BsgEvnXCeDSF1vrESiV
faN0+g6iGn68j/u4D5n9/Kjcl/XhizIDN8PtMixIJgl9AajZfx8dSHFzrZ44CUXWyEsdnyVp1jeu
GXEvfFgkhSFTZVbdDTs9q7bHaK+fT6O+XErVN6CW6UHpuSFsuBS09keGdZ6lipN45Uj0yXisNYoy
mf2mXshJYwpkjiu+NbziGQ3/uQcIzIz/sZUQvGo+ivZSevwR25Vd9HX8YWRmspomRaOdfPQGAg/r
rQZ0YE3MHeiXgqOaA2llDn8v7I9pKMqerg5x270zCSl8BogohiQEfk3qvnJzP5uoY7Y/I9TPfs3O
aV46TJDKqNTfn0zgF4BpDAFBBeR0Zykf+qtDXVGfYhrtquy4q2AI4QF1KaoYiotBoFS5Qm+UyzWl
VCwYvT3WPXZFJcUMdfSedVn7TLSCornbkiEjWRZ7FgdNG1Do8kgeZiQK7b0dYXp+PIQnyi5JrgCa
MRlRxjjtUnivG+ajKzo6UpKxThVfYuwJwc/58JGqgq73XxSh+i3vQtGEm67FfMWpy+JeIzms1nVm
c2w3zys9jEchAQ2iUoG1k8w2SmMVePH2DftrJg65nY4u64pvicpECQD7jR4fF+w44zUFL7WXnp+b
Xw5TZJrbpeiQcxpPCbYXxrb2Ir6zWNff+LGdfu58SLNsKpLL8IMxMDkdN52/S54S3rXptNOad/Rh
iAev9n3I7Unm61kpuOo0Tu1HmerdwxQJIdTtDkJgFsF6y8Ltx/kQybQv2BD7cONCqIAF7aowEx1W
fl/26Rise6poksvOi63TwIIWRLnVJJMlUKRpeTc7OFdpRCdiDMWt4UQfFxnXDZ0+X6BG9HPyErtf
xhkIuTouP09zoQytHoyAE/TtCFBf8V7p12X8U4oMjXHDIloArwlWeySv4VFsdt4HKfXHHm/5OkXt
C7AHvOCCcJlyKet1hINPpgWPJrcrp3HZPn73KlSAiLJsMEDM8L5NDOgyzAH6KSsiyl4DfVL3nlcT
ramiLInLDBRdxw8JwDZ75A7z1XPE1J0IUtTWMhwgvGPOgY1fLVJgmHDSYcDD63QzUKbl5OOALIWy
uc/bWuzHujS/Enaj4jnWEEIllIgR3q4t2kutZTI5L4Q0Q+3jcIWaSOToT7NBphf7FB6baz+CpWRu
4YOPiV8obs0mWpERVPPkFH3hmf7LkpTb0TJGoCgSykKCO3LztJQ9KUlXFXWV0UCeyj3ocryVfVxB
qXaBvwVvBnSsvSiwWOvEXfDWF9rdHr6tNc6BKEWtgskXLPopOPhCBF1fmzMvPJK+Zr5WyL+fmMun
NF/veNw8W4gHBFuJ07ulQ0BtuV/ruS3XVtJ8J/EjBQGW+wVpSJMAR14zbkkr4tOpKkpJ50MySKyo
WfIZMXNfAEjdpMGQKv3B8CBOXtUcZBuwVJeYrKEnrXRl5yHq5o0+aSwTMcyWmfXDKUhmkESksuho
sS8+NO4eI6BFh5Smz6hLDjQJzFVcHLIckZleYdMigxFDVp0art2W2hTsseLcreGqGxwzjpHbeXY5
pYdqGGo1qipSyOQmg/RHbtS7fO5CPlXmr4MBGH7HwJFYR0OTS5iYApBzvjndvZ9fCoNtkLDQy8Bo
5JMtrjZIuN6uMXljPddPOT9RFFVw5+NSp2v74DRPVU5N8gGBMfCQT173l9Dnr8dc/nGsBwQA2/eX
qY0zZ3rz7ULTGcwz7NbA0rhDKUHw0JwAv511Nw46F1/wXE689hayWQrzan7gWhGzEj/0HsmlLoDd
96J1t1mQpRCnF0rfKbiRMgiie6v9CjLY7uLNtno1BdwinjN62F7091xCXALV04UhedFFmFPUgjzD
yK2JCE0v0Xky5WsmgXd+38m6fnb/bmVjHf/lXH9gKoKj6enRYGzPHyjir/sFVeLqeiGoLIn9bL2j
vA09/GiF+SUKlDjHlLT3iQh6sHSAG8Wh+uqG3p84b8ktiTmtNm0ASNf79i2ntc1L2SViBDibWWG1
NmvD+MxKR2lILAj5QCwVyavktnyyPGIocWOOKzYyyRTsD2HBOaJDjkaMy05A5+nxHThapV+b2oz4
QcSbI8PDH2vim18ElqFzn41+mvMYk7Rure1er4VGS39z4VRdit9NS9IJDPItTwWUBL7QoQX+hvJj
Q4T8B4amjoZiq5YQjfPFABkL7GXgXAJZavZt6ecjaqdQO48ZY7zgl60ehfOyXuv/NFNMeweSjHSB
V/CdwM+f1jCwwRv6JG9Lx9ULRhfAc5ec4mYKqes+Q+kv5YbgJGo9YzmniyowDThDnxtnpEd3l6yO
Vl6nlO1fkEO9CuO/8WeTLiRgYO1691VoAfSstAiaDDFnE6zyCTycGg1Gg5vOe3mX0Gs07jeQrYMp
kShFIHsnnk1jFQL6Vwua1G8O89QuGwIzHYzx/SZ7AsvkT20vzmJORMVyB2wL8KQ1tdO3JT/kKaf0
PPngk7RXp8u+YgwCqQ8PxEhrWICS78kUNQDzsrv3OeUR7UZOnhvU+QttWa+f+ZTKj2ROWsfxIeHW
jbHm51BiLfIp3+9wrLAAZBB2lyVw8ZC1p13SmzJzH76Mml713oRCadEdymZtd23DtS3D77pzCY1S
jzOs8OJDE+346BlkoPosAmpYizKOi4mzAWyKfpDBbE9PGNXGePVhJQ5eAKRWrGBRedOK5etsjnmY
LfX9Kuhv2imCCimVNQkL7gsTI4JSdnN+R9Iy5W2RXwXS7jFws8YktI2ttnt2dwgxbCkCBWl6h9Wg
f1l2R/T/wMe7e6fkmKRCggl4XSmsvHzOoy/8FuWARdvss1fPJe9moX7i4t1eUK7xVgCF+7RWnmWJ
Pl+KDFXPwis4rPzPRyiVwZKnA3RV+GlgK/XqIEEGb9fRjTL7jsscEDlo06XeqSnADyx1rG8IsaGT
bRby5vGrEStT/YamYW+Zrv75y3lnVtUrjMTjSVatx577/4tLSMrowHTC6/MzC/ya5MQvt7CHJIBF
V8fW1b7zOp08obCnjwc4RhXSA88sGEVjrH1ShjgvUHJkgZ2mZ56NrVX7obg6I/AWXHLzZ+p46GrB
WqNCJqsT9a3eMFl/ZZnMD5oUjYbaCIgbPUNLhkFQIlnu374Z+yBPmTIBtbooLApZ53ZIpEk8R1FY
nIEa2V7g/WkryObBchdF6r6NSVr8K3kiU/zlxmzrbgFc+RW7OHNWjHCrh2CwOqLfhajMopxkZa0a
F8ko+mUbC+docObLEDhDCis1jp+zAVzCbJtveiHqf1xxw+rE+jx0pjtVu+v0CInfQdHsl8DxevN8
TGZX9m/EG+cWkrGNXDH+ysmhGJFFQ89eSIpQWrhpTfO3831zglGhmBuzHMByRyx5QypkJc+pZYIY
GNmTjdJo3InkUjk3CObTV3Uez8lgj4d77OQ3/1AsVV2Xlvoi3AQ+0IGnY0K5w22cyaImjWPg8LmP
iHgmcimOgRsc2KI8y9/Hb1eVl7KM6urA1svhC5BeWx3CSoXYGb6q1qoHV/+ZyB1EKWtEuxmcitzz
H2tCB/81QzWdaAyMu2koGyzeTg5CIRnMdvOvcZZHBvuT2qYtcS6OJd1CgPkaQOmP6ySoMJv2z/uq
ubQa1QAPgLuMYyzHMBVDm5hqRy0g222ApK/DNw6/NUVfl305y0rA1y73PfxWbD1C4sqeltrPP2JQ
pUjvv1nlhoL6i8+GSnOykoTq4dFi2Pag3uz9Ol9ezhNvItSFKCRgAMa8fMUIKyQJnXsAdY1sAWDY
/HpoKwwmk/OXG/JWr4AQ6Z2hz+cNyD9JEiSc6ENkZVxEu0amRO/oaNHx4GciPH2osTkM8g4eyevt
dLlMF8fWHlZJT3LfN9YaFaZwUAWFDGeKdfDwpl/WxRa7zqjNiGDY/iCImM+yfXDDxc4Xi56l6RK4
gkLZ5Ln33R3tqo64e5CKjmYKc1WVifr2kH0I99f29MNxRwv3DGYYWlbehGQZpw2a9zMMfA9lo8nK
iJbhCH66vrlWKJgnJxmQClSoyOKOQG8gE0lpcfEhm1CNZWUYl5n0iL3ZjL0pC78/GjpCfVIbnXhl
/nEdP7ELyKV7NftWXPQdGCba2RH4TrSdaOFOg6ArAX0+IrO3r8KkQotOTyDnrMqfjc7qYlA4O1KK
GzQX77KCEmx4XSIzYrM7AgtMm1o0aMEwwwH5gzfRVhcy+Hzwrox5hkvXBSt2Pa7W2A6UuwaeJKvy
6EzrBLZnNic+SDjqjbItiuCd3nilJmqd8a0zO8n+IJ9UZ3OM4GsVM4WWOXYMZBgaf8KN+vgKUSDM
2MzvXaR1Klf7JakgoWkdBNWiPPiskxNK5omL3ZdJ+8vd8Iy/d9LDB6HIlTSQ0QR0DAjImhBDNPaK
/e0OyfriMQrMjctsIXHKygr/8aXUcK2a5Use/eyFfniFQ/VsaXM8Zgz0kzy7ooBZMckw+qU6HFKu
xAkHb72PmXOwnp8ddM42O/6AYRPwWyzt9KW2+xeoOywswWz275qfKIqOayQePnryvTquG3ok3yI8
rLhdDIrfFGrTnLdS/oDx5XDENC8aCWcRBhVzvb+9FAjzzpmVJniH2KPFj5VrBkVrJGOKkSslK0w2
3m9S5XJjjb5vMOOh7mfjDLqMZJA0G05S735Cv92JvpQvzU2uuCQqTGmZ2OE6PV8svsj9O0GkCE1o
+uwkD2DV/32HpjDO4PUAZ29zrvT+RZiPWtJ8Lge5aadiE1IV/BZSGfoC0nzIRzytCw7Cm1ez4OWC
chNELoDUOK2Raoi0iZ9OZLI+0ABgoJgokfsh5f8PPoUh5CKtcluA/TqN5mCCGQLXP51mpIdWYYNB
Rte2QznCwqggAqx2+gJW5XczVGldnQgCTYyazGwrfyR35K3fzWWUpNsnMx6M+nnzHMtcK84TrKIq
a+QglpZKWuNHtiQ4cwRCxoM42aNnYhj5vaZl3i7HgrCdwz973+rVviiFM7VSqvm/cSICVtcp3GKL
Rxc8QxW9mryNo+EOLwZi20tG2zr7bmmpaV3avm5JOF8Ae9uUI00oka3Jexe3zyzr0czwmW+NvL4k
NHR4xvz0FYzOcJdfTG9KfZsJloPFTe0C6sw8w83FXWFkUIt822orUxyQPEWBc1VUFOOx9jQrezSu
OomYo23soJuUhfbLa5EUxDZTItocfmPqaRF07Kfe2c762H6rnUHVZSKGRxWlRksn/ddwP30gIziQ
cXDOvwNt7O7etYVNXrATB/FEn1rmixn6x88KZYlzzimGyv6hfBorkxR1xJP2IEJl7d2BA3RRW1KT
ZvF2WqhjeavkFPVZGxS+kPh8eYBSjvV7E8hcRy5HitHMzZrBZNC0IWK2IBLB4wfnfCvmf+BxarOt
WteBtXXGy+7/fCgiZItGfMDSOtSAqI0g/ZdylfC4ZnxzFNmB492jza5I5cIDkjhDuvD3lWv8edg3
z8KzZB2Y4iboQSNh/3YP36M/6xQg701rqzX2Cmf1TufPkUuhjGOmNWjq3D8yBsXJkLKN0zPTEeym
qsQ1AnIJkKOx+6UokUahLOn/uZkL6GqIBHmF6d3+NuINKzUyPAJBZlvoevTzTas61/g4o83v9eRC
j2GsGX4g/AEJTAdI1GbP0jFjnjrCyx7hiMzqQqp98SYwdkUCFp7lVphCoMcAhFUl1DpmV2x6Zy9/
gWxk7JWwSs3xsoRmis1rvFxuGF9ABWG2MxftiOtPAgmDV7dcLHkKpWcq47heDdF10xQIAUWJQhJv
CBQ4WJ0QU7D7e7ctzlIjtlInb7P6N/79/ZZvH6lnLUER6nvEcM12+sSoeDC7pn7OPr6pIp6En9nP
HXcS2TfUWzHnF7eK7YBGkQOH0S8WH3rEhb+eynNM4zTHdSsqIdJxJKKlG6LNbeZ7WkqY/45QZvTI
yC1+xul7MQ8ReneM9aK0STjsHRcP+IQPigDEBJWCsyc2uvPTuEX9ZPxdtR/iItbr5u8TbbmYSKBv
aFi2IRWH8pcubx93VxlXhF25rv5UxQKrqs/cKrDFPk2nbSwfo5csbium6RaQr5T4x3El0p6fs6Oj
+dpXsMaC2+8PAtmhkSUybzUIWz/kuHcXvd0tqVrmb75HVownyyRly+92mWoc+Te/dUqll6pTp1S7
rOPEEgUapeFCFFKinCLQ4bD687qzdjx3bD//yCAPny4wfbKJnnAlq9CQjkCymGseYepfnCqmcbfJ
TIQlseQ24xZrGjfp+491owNJ+UUzRW6zLSngAfX5gkRmVKfvRAIRxrOTv7a5ODIv1YAZRFjNPX8V
2MD8istqMQRC4nN+w4d1X67B88I5WnY2v2YSFORhwYhvueB3muiVmSN05jOrQVLjJiPrXVCweEy/
sZwyIn8Ka2wE0uqqL+mW/pMmo1gzdzT0t+Gxz/t89fTzrzKjbIUbLe9KUEPWGwQKDjeGPCUGvLmQ
DVZR2YUG0yhcttSGFtvFffGLzubp8bAC/jhIzW2O4katXBpfEor0mmhdXerVvVTe3t5rR/tsN/hS
nNWnjfjOOhIbyuokflpicyMR5n0j7mixS1Z7wizHjXY14xWwLDuz9YBtr3boWZdXrQoXzol4qUJO
n4k++otzwYRIrNVxYc3OeNOzHueA5sX0do1HECA/DRMMIal4oOHQlSQMAkCpTkJTFpy4LN08Ir4W
cvYtip/B1/twLH3nCb9wGR6sqx4qOdLsw2I0PtzDO3lAC7xIk31ZwIoIPc0S3Vmq8jzm8D2O5wqE
Uqh60WBlbrJYutPfG8b3SMKajn4Zg1rwoyuXObm0KlFeixNrzK2pO+nlUZt7GQ8wBeZBMEM63M61
hYigvNGFzSzNcWjAEOMznWoHqSNkl2kS+kvAFUoyYDYLOYGDXvB7Zq5vxDGB7Yjh1w7s9Uydl+y8
ScQqAPhBiqPOYULZEkXOX/jkrxf7dX9rRICHDXHu/yl1Wdk89P3AMheOz2L44gtXmQrLOb2ZxHlR
s/pYyVRUKfqgga6LzMJOwHOp+e5Fn1hs4eaSDLaV3MvIfXRPP9luEvc7Nb4qy6o21AtzLPGW2djE
t+llU1bQ64YESGn7LHVrODDW5pLYI/TC8Kl4tcWavMTUu0arx30KUKTSH4wPUZnQKdzEDdViZ2Ah
gS5+3biJVcPlBz43LelcGl7egPpoxRC1+VqmFd/yXEZAEPbvXudvmVugvYFHpjuX7h4iaI0CBAw1
Er3HLD3eSpPT5wf5VhUmh65YA3jiol1/fApnoNe2UC+DZE9f+4E2ryhJt98enQg1V7WHXXZ6ZVFj
z+jjpUP9PRwJn5oiZ260KxJuA9a9NFAR9/JRTuaI/gtlYWtC/l4mGQo3yMfZbZCumlJCK56xATpm
OLiE09Ryl0rVbc/a73XzYqn+PZzz2bK6FhiP+144wbMh2Z2UnoNyytGafZconnQVD67F/SKvVnnQ
xTJ4cmNEquJ5jeMsPiHLRbijfuCnHfZhB+fRPtNMLyRDYhgD6cH/KJpc/6W1kSllA7+/4Yef0gka
tPjgHKZU58c4XTKM2civfIKqR3DotZ1YO1OGRwRqXMkKbnMSqwWyo0tXk8OgIubKowu7beAFBnfK
JzLCHYZGzlMi2BVq86mYWz6y/vJoLslf+xyVK3E1FX+sYaaCujHfDSHmYa/jBjugmAQaOE5urvsM
mRXSofNXmYHLza6RkznjLjukZKBiuut4jGXzma0eUsCcLeult8+yYS+Sza/4b8pE4Ggib8tVcUud
COckY/LGyS7wDt5RR/6ggovp3edTnV12ae3eJyOBSuoTMiJkxfjbdVWmdxuBaffJMbo3UozWzTT4
SJNLmR00xWplo/gawmS8XB8ibpcvp4SJWGrwwJqot5XVZM930ejLRv+zV4vV6+Tv0muX38Zh6mRQ
XKIrLC00VONL69ignPRln2XbspDMELqhq91Kv9KPkvOszLYSm5GUBQZ0GohnIBSVMSTzTWvaa7/A
kyw7p/0LDu01am9aC4O8kne2XWLgJuelrnCFtsFXJJQ+zuHZ7uD592E3qYAKhRbb1BBE5lu2Es7a
J6QjFtQVKbhgjKpDQMVER35z3bk50vYn8Rscs585BVffcSA+PaRkdQFYyVz3smM3WV3gRTOYMMLA
DI8GaeOvGrGjCO/jdruv2kCHBb4FDEfbdE56icjEbjMMwfkQ4YbIX17avh2jKdGSuj4Pz2kP0Ir9
jwlyQPrOKCm9hIy/VEVZoDogCdjEW2BfwIWFZ+SXosQTab6MVq5UdWpPfNzPUwJJ1kfghMBPv53b
WwJBervzXX+EX0ysqf9mGmasfTWY31siUtPqExrnC3MeSbBwOuY9m56rfDJ0uGt1et7VOr2Ro7Dk
o04ur+2Bld4w4fdpaiktKAnSCT7W18nihcoREkMn7xnAWCIa8VRWSd+jTOI2k+AY853SW8aaU/z1
jcsMtRZCN81eKkgqhCvxPmvQ3bNLP2aABL+GkmCpRza+H8npMoinqg+OML6N20bcqWt8gtilOfdr
Klj0kbrM1cGavdXb7vx4voEQEpP7ODWi/UQthXc1RO6OGNL/+2RVP5veJhDYhllIZoWiWuS8y0XC
6UxyfjwT5TF88cuEpQTKCjVAS/C844StI4JsLYxb7MZwJlKV6y+WHqYuznEfTQvMdZVa4xhrvLBF
8bJ4/0AX0XnzdUS69TX9u1Ifn5PPLbq4NSCHk//jjiX19942iZKhBrTQKD64p6AoXqgczTF+XbdE
Y81uiST8G1bGNOVnZBUO+rrQsz9GJ4QC2OlAP2tHLoDCsplXs7vyxCNb4msogb48eXO1pb98E8Ti
8O/urqABr7XgEw42FEYRy8Z4Vb3U09Hg5emboHejzXy3ebpjZlXobc7XwG2HVvYKHdeAbj/oewbn
78O2NjLdHjl+HPeZPGE0YpOzLc5fJinnAGYlASjwlVz7PJ3vZu5QKKY4aOyGZd+f6v9hxTsW+sWh
jXLrwewFrGriMuqMc2TyDAxm36bPqE2mxDWqzUiTptAoKjNFyS6fiY6Q8HbTtaRhqgaaRepsaI7b
VQnTzpXqCJUkoboA647IddpaDxjNTmL0F/OpAicJ1fqNxdo7iJoSF01FBY48gck95BKDeR/Siey2
BAFJrYUoc3PiJ+jsLgSS49uf2ixTGFh5YYVmRMlaBvhpFRbQi037mRM4EdwA4jL5BLDBh4XJoqSO
/hXk6yGjKVbDaQAgXz8eNHdI6sowArXte36s5QWxQJF1GOR5SQPtcjY2JcgI1fdXyoLQGL0XuQOA
GywodAMYMgCRG6KaQ1+igc14jeHeGwSBErmLd87FhfWfWJGHgEiCZJANK/uqY2ykgdEbe8JodRmA
LjKa7k34+qQOkOBSxU/el7ddHfl4c8pzLqbOEhOtQJ/6ly8EXrIIjYeyjsIGPZL5CSOHzCBbFtoZ
HyjH3XmLA80RFAzrh/M2EpvjQi8xhuxU6HuMXWIxP6lYqn1DN1oByqLxkSlZEwRcVVlhE645/qeH
Oli93lTWfyo0cLBaijuWRO2najBLvyyFzTJBM9w5dqt4t5dpHqqUK4onUra77G0T2+QZSuSBcaCc
MX24snwHKf5Dzk2gKisANMZzzyMsuR4x7xd2Bc4ru9I63WAUtJoA8elJ4pqdmPiZK6iahXttvvH3
NBDEyWzbepVjUXHP2hbiRcTdHLPLmM+f1ULDcuRStwBgNCgS908ZlWevAU5gqscroMri5GYMcFs9
G60H1QFTWEyOaDFCpj6mG5deCKfAgBYSA1HgjXlZUi5f0fRWaX+nb8/sHJcZNT/GQDhNJ4m9XqSp
SfUwCHQRwkoYkvHzWriHlTmHdG33Gpr5NYPrCteGU9VE7WSVrT4QKUwEttSFENtSIUyVuSlqXCQV
Do3NDPK98Z1yKZ8xAh6ASwm56hP8Kg4aWUahhOrevArnfE6X8txdLOBac4zeJm3lUtF14aUPznOD
ADhpvhr+s0ZbQmpUntVprJTubT6oh4ul9cMuL7BJ1LiM2mhdxJy/jCH8qNjUhUCRBkCVdPA5r9T7
2hzReBApl5hjDdEPv/UMBMRGr0d4IzXmQstxsW+rjFMhSZkZE7Q+dxrGO3XmHMSFH7Cb4E3sflen
fv3vxLXPV+9Ude0hG/MrHbpIkocrVqEDWmsuPtP9cwWWOisLwRj+KVd5wpm3Va2iyimIwO8a1d3f
9rELpp8ae9CsBP7fJDH4KWS/SlkgspGgsR9SL5Ri2vQszM0RpzpvojD13JaHyGkLYculnKoRH2v/
I9ryb+K70JaYu+awMpzvl5O2rfe8wau+jZ4HJzy3+Qe4+d5SZ0tMe2FqMFPTB3C4yyM4hUZMpLgK
Vdzy/gOSqrpXVQ0qSlY4fmvBaY3/gcyej+FrsL2hxz9Wox8SC2s+5mTt1EBhDh9NUS8QvAPzJ5MB
14P6rBkgYMOv/3W/ZQvHFcW9Jn5guUguTAB0zDX26dOFR/KSx7M2+KWEPSOhulLgUD90+kYIHa9R
A9z7rwpgvMeEn0DH6xCXNgDpotJFswdsVeO+yABH/B5K0xFONXaTGqm/ySJQmFd3JNnQb+3njy3J
PaBe3D7seQnKYL94zROF68ueDiFJ0zwj4mkBNJAqMKpMvzo9r5+5NtgOuxMBYX4iP8/8a34C1DIN
QQRqrOE55ZlJ0wEkueflnLj3tDEfJMnDW6YsqlKFXzL58gsgupNdzhMUWJCkWlUFYBOb7EdvCDM8
yqmCnxHH1XFMZLwNzTPVKDdfIOelJxp3IKTRnjlG4Qu4/xm4LfI7/QiPt3aZKXWGfAvyjndJFcBL
2vvJv2tTC56RM8cPrlE1QMPzEOpccF+lNz59r0yfF0Jx0zA+DxKAMTa+1ld273KOcNSsx0hpi4aq
q8aGUA6RoxGDwXBD2Rea5T9pMs95R9HrG93ZQhZ/Akbdtnry1IkTwTAyw/qd74gLkgRT1lWDRkPj
f1VJ7Mhxf033jSnScYIGzx7uRA0o+Mer8OyGlcmQYlU9pfWD3xfYdXdujriNQlJMT9WEcE3ZEm5c
7RHSthqOFeT0NSaLoFMiP5d6kfu4Kdc8DSLNCisK8EoiH9oGrwzYaXwRtrvDkzDgSxBgVDA4Ags0
y3lu1o05Xbs9tz7gb3Zp0PT4WjVi0/ca8oaobpkMpiJFrA1jVxngrN8NjYjXxmb6bIdiJN/CQTdX
Pqwpoa3ewB85s7jRVUzgFkgPC/sMnUQEfWePVWape9oVkZGDeexS/GrTeF60kDUZCs2pFMbCQzwW
M3oeUT2nhP9XwuWtIwrThubE/jI2O6mQZWD/+6L/mm1ni/wbkUT0DvCFFLQYpFvupYAIBwRgfrcA
bW1NOYL8S7u8R2xr+5D2eDd0j0/NsYNf+gH2GxjyTQXhWnO1S13HchSfD4aHpadCVRPbINAW9IJL
oPmGTe+bGHe0cAL3XNMar7tXXYJS6f4jumQBUmyRtoHNrA6BVuYRqUOO7BZHRMM+WtstGwbjt9kC
7ObA9OQNwV/Xd70Sfaxydki7DluDH2tECuGdxF2dvauZ/ZF7Az86DIM4daQ29qsKorgIqYYxZkQf
U4K8QRziH7C6DuC7O/e3JHuuTGAP2ddyhMy5368hmMSa/hQKSEKqN6wHr4aWrca4wcQLjYD4WSNE
GYi2t/GJBoB5DbiQ2gczDFaxgFCBHlsBDSDoIu0MxqqfMEkmMrbN2WVtOFSu2R4aDRLelRjUVX8k
1u0F3KwNlLIq5nm8qgM3/UtCc4bwhguPM3pqYoF6nBNM+Xsu4OcfmU4cll9OvdP59I91KRtqrCSq
rD6q49KTatBEessOmax6eVJyN4Pjs84j7ZbBb5w/NXW9531HtJmFGqVF3oeWVFTjvKgc1LjJIrrb
w3Ulo/trqkObQeTXivbjHFABx8elo3fk3PQ36m+AYBrRMydiWOhVoeTaGSz1j6bf7v05MR38MrPh
1d8bpZqB/u1kAglReQrERY5lgDzhyzjfsQQEHAYQIC3xopHpRn5VouGnTEPsNXB8PaBiuHTu0auy
lj6MML2qkAITBz9O+YQqKpEMMgliSBOtOxW2387TGfnF1Tc3znUX23L2dECPfvEMf6TquYH0ovW1
2Wxy8TVMtfEuZ6aS6jg7t4CciQCeoIgOWusJdC4GLFPc+pz9Je9zZYvwn38lYPKPgRDzJlEvGdbt
sYZeREzn53qUN54Z4R8y3l7iEFjgu0OmKuGN0F5B64HWyuzEy1i2mY1O6a2kyZF7za95d0gETr+9
iWqNCyi5eHZKo8YYJM+Oc6j0yzh6ttmDtqr/VTlgbh+zFGBJMfsb53tR3pBKXIy4V18zsj9uHz8b
DVeQ4Sc6rSjC/N2EipPuF69fi4/Y8TCtMxfe7dCjv0bTWrw2c/o+uVVl+WbThNDf+4vkprinXkrr
TyFaW0kM1vjeb52RruPckgjV/xMJqtKlaHxgcKYOYK0c2WTr92UT7XIZft8h1aYPy4kVIkvh7GmX
Jr3txN4uJM0+6ASPlWSaxIR2bb4F5/bVxV0KFKv391+73d/wMStJKUNq3N03XsfYxAQdYz7V13XU
G5vSTkJQGXIRj+Dqe9/ig5AeWGlgnwYMHq3lYxIUulFx/kLnOU6DUo3D1t16UcMvG8w0y0bDkFvS
ghLMIpyH9SOZ5sedyseHV/7CT+Hy3iH9iWElgYbks0gUcK9kDiP+ZUbhdrpLrWuzmfXfgQQrmrqj
mVV7GMM4Au8akABw4hbuYNlJ9hqFwZfpHPXtI8YfdMnVnRxvkyn5yAoxg/UkHdtI3JB1oYRKtZgw
/RO2ZTPjZ+bJVeszX5rkrGMIueRSFJGVMZPg/QhegOBhaOeIxmjKctcBO/+bd70neCn47YabDvLw
nvR85LgPmFXhd46RCqAQnOvBK6lWaRzN9ud3HFXkVL8K8X45pFFwF4Opt5rZcyNajyRlB7X1+MKK
tFRIhzyPHYlYabImLYtprNI7N6Sn0cVDb5s7IE9JSq+aUHZfPYMxjO6tz1u8bPT68xqMdFk2ZLBE
9ApPPrjODDl+MIU4wKDQ74lhaEDxFfo9u2kpN4jyg0+ZVavWf8q7/p5FNzM8sSIUdAU6o7QT9I3W
Sb1QY4JbsQNXWaSP9augajLQxQa4Knw4r/JBpB+JRObHxfbD/Gztf3+zMekzDEcq5bfwWeT5uYap
teaX3kPD2VTellzme5GwC0qijNzd+QYJtcsZoNdxl5CuCHQWrHCXSJjX9y9eoeoLUUxTPjNSJxIx
aP/WefOrj5U1ZlgHQQZOBYRaK/9O1G7mleibqCly4MMkNWpNjzmmxe1pM3uQ23f2klPBAeZmiOpH
ZOMMZ/LGYg4PlnvGGTwNuWlijeVGP3xgsyo8XMmPI+Y1FiykdZYuID2BScq4RfMPi2XrxdAyhjie
Ns52HqQuedhB32mcr9cT/SJ6DL/wbD9F9r2RdJ/T58oleOwfJF5eOA1GcW9XebqUCo31Ky3XG1XR
8BsYVutoR3infRrSglcs4v3BuovVt8MnFJPQ7JjLxjxFl4dk+HEVIaf+ots6HDItsurfTA3qBZun
qD1xZ2VPlq6Px9DdKHOXWXcrW8dKLpO5v/W18TIw5e1hfh5IZY00LyH6sMhTH4Ef+x172qCsRsW4
kwvVbZcGz9MUEdTb67Rs32uoDH+pAnArPfdnQ6UbEzGcqXsMOBYGvJP8jZRPbZRAGWvir7JAnD33
tAhEZ3u3hVSmKaEO28RMK/jrJ5B6kxqZzgnFUVKbuhIf47idOzHq69LihZQUHn+d8P1dT2cfu7gr
3n1M8mgJcxS6Yy/Lv/x0w3Xt3DZ/s+0x0Vrfr7lfodYpLPcZNI30m61nYp5/7sscm4BRBaYloexN
JqpNDFKldU+2hhGejPowFis/kHPjgn+IZgdFdkilXxZuAZlWJxj1p3mNEf1fbfYf4r9azBssQLAw
TH2KoB/8H4T2FVMcxdVF6WXph2aIGze9nv0poUzZO38eHMgsrHazJ7H+0Q2GdfBGXredGs77FotA
L8MGIptFtGn+AiCmf1dxNgsC8xSWocOixrZmf97dyxlO2dB0aFPQY7vrrd8f91xwGy9seAsbiuLL
oa3VspGxzBrs6e6+RiM0d3yu5028Q1OCF8EBScYFrGftwasX0sz/WODIJrKrtTwqwbEaS1Jbbi4q
WECjQB3xmmd97EQKGlpKbriCGjZVWDv2NKGVH1xbuV2fh+eAjaT9eHdauPuZahPtw4xZ0Mpwk/SV
zHxg3zXY3Ip/AiQ7zfuKpsBuBOqXIHY1+5SZhFB2OYgu/hoBQ0OZ7kbF75czjQlBOYqpRJE57N6G
MzlpAP/3sttx30gS/F/vOQbgp9lVjbOH+FLOo9m5k7ktXXyhxbIOF7WStajTe/2zyumYldIv8yjK
ZHqy5sEGxJyyX6oM//CJYu3hQZU+IzJjvbRLzRSEu7QcgWoImtdh973UQ4OXRu3I+shORFvDM9uk
R6mClv+9FKwMGeAFabLk8lpajjbQELUakkZfqKGnHu4TVtL07G2Q9RcF3rFmd07NFFeWxeBKg8I0
MW2HvROiwIEZQQQntQbjen8Sh5xtKB/oTGRDS4mCWVJl8y3Z6rNyPTnEnaSPCTmhop0noSWbZWLg
fC8l8iCv5IiH94+A8VB/9wyvlFEJyQu6LPsEVd7r638Vh03ieKcZL1fa6MWNY1rFVB4aNR6Fddlr
MoWS3klNJVg0TrtIqHMcWOv33T9o+yTQs+nsQ2zLKW4d5Ix3I6D/U3dwPgKTQ6K3K2nhaQ9bGoCV
PwUEvZP/6p/g9oAAxRTv75tNnSo6opBLrOth8IObGJQNvTQ+3kEI3pdNzjGFbkbKsiAV6RZXGvEe
nHPjJEYgU4B2jJ/4daoSiDerJEiESxAb+yA9+CXzvcAW1DS63msCiA9oOSCaGj/bJiluvDCQrh7J
N6OluVE+W6bIY/EEGCFyt9drGfKVa6SleghAo2H3owrKD4jjDuqd4W614ZPhpBdOwzu+D/sczOO/
6vyM2Cugws+Ir8IpHocCzPGVSpgF7ll0NQcjFY6dKvkKccspYrtHKWgyTtteb+SLbU2Sbvx+tDnF
VUGCaB6VScdNU9JHJK9jiE/i9PSJo8ddqnidNJv0DK1H//bPlG2Nqpxw+AGDAFgNMmdPxqVpzZ9n
JCd2k3dz68nR5eemBMbTEhl2EI+2E3Gm8D5/xTh9S6nzzfvwwxJcp1robwZdya3XyqVVv45tFlFZ
lGqcNIix7c4BLYx2JVUqqxSJHURIRg/0r/MclIbUhNWIK/J6YuobPje0VP2Qh5SdIQx20FTowZLX
2giURrLPiN9O1dq+ekrSL1ZZqV5vNXa5z9V6ssLTvYBO2GKxAnzk4HjTISx290m0GwTDGAH/3xiA
N1DmogD7M+EbjFFmkE1zGeWWPWn2lVcEFcDhR+XUIdlhAEur1cPO1LJnSEpoN9iGGM9HiQboR0pA
oLNmN3dr5X+U7pC+/ieIfFoRleXY/2OslmCXtevmYEuYGITpQQZ+ToXF3QLMg64Z/eY5S1xg/PFb
W/B8PTZ51j5gbSkQVI6JTSJ6hl1Y5nQk65PObx+gCfANs+f6qywYpk79YHKcdg3burmbhLTU82BW
3UCgmwhKL6kA1zFDgwUWHrjRT+5leDw9TuCskpaYNqruAKFwBq0IiGIyQ90RjtXMB2LUsVz4XJIt
Ki1/LfHMlaob58nYABKIuow//MiFzKQ/lQF6GTz6nchwppmpoDXN3mPRzlOjtK4OxuhYF0p80mkN
R0pQrRy91XHpma933I77RaTzdL+7MMKw4SUVsMfSP49iZTwS9mu/zimGs7V5ZxvFahSYrD+elHJJ
UkIWVTnalaga2+53gh9tA0nFk9ZueXBjw5ecY1PWwNGPtRJb4zcHlx9igas4ee9zuv/Kqnn0CP2L
Pl25EdR4vGVDpeuq2hSA8FB9KQi0r2hrBjotlYENSHX3hLhHpaVQIYuOMxzfMoFYRnFjKcUS3OCv
zjJk90Kbqn28B+7smKR/C+iDTDDUV8YVKSLqaipKfx8eZYcPF6ZgI0VwYv83RurxUCjNCY7eCxAD
uOQ9bn2/DvIoAFXecDi4fbbbYz6Uf3fPpLTLnAQmDrLQW4OQ9mL/dEyXjqpGgKpXOwSy0lXDQRoW
vW/7rSsNk43LTvjHzXVcQ3Z3uZe6x+uxt+2DO4S/QgEMYtA6M1k+1FeCQvHZS72aUvWRgBW2AE8f
tQcRl1YIQdLD7RLZYJd+gYNYeu6Haa5bvZpXDO2IbH1XSBfooM8mefar221/kQPTDigqqivcDH/H
7M1KkYcg+KRhFCjR4JdCny6Va2QnlQD+ANijOHraT5hUJHlamTX26ipEXpD5JcYQdI2xAUNTjRaV
WEqeItukzwdnQGtRurV9t2ZEQF6kuYlyD/SCYW9otobQG8dkyTJMMpw5fmzAldI3ymBT0pYNEs42
4U/82Yc4MbHW5EPNNNlgMQyuPGCKIZZu4BU5bdWyOjjEsEiXolztAEIRxqA6R65YAyVmO/xSaiUU
ho0hyJL7DXs0ofGDj8Nn9w0yZ7Q/mcvci9mxrAKu/T8NCZ4MlyqlcCpP5B9qgPN/BNan47zvMXlu
h81wyi3pohf8i6Fl/2jcMsfacqSj8ADW33LedhVclxQBsdBOayIFdGYLwNkWSl3I01uHkZcANWGk
V16Mbs1YOgTxy4nbHM2OGazxZliuZucdlVWtscbn3DxybgMUZ5jgwffqLRaRWmVV2jrH4FNciYVl
fCLx2o9gm/zMQighukvCaXpfWlcrRfugiEnCSB5B2SFzSltHxUmz16xSewRja4Gwb2tp4sj/BVvW
VqZfSArYDP240hhYutDQdWfIwFb2JyuI2J3xeMR/28PT+iiSWjkU08/w86dP04biXEDXPS11wyvC
zJuefZMUjKfYq37++8m+LGomFEVqnZ5HTEFXd5VjXrQqM54hNnraTCPqOGRzSoGTOia/4PIxe408
mgO/w8KuF66Fk7NRxduU8c5mLL8IoOXjBNUKX22hPYPYl1mAwJgQQAE2Qsg6D0RMwF7quW0foY83
BKLb5Y7PXTusf6LvJ2n6AFaPs5YBZZ2CANgxgIlYkmYpHhIoLA1iT74tta6Epq3j5/nn3G+3R71u
5YwmhDpfoLPqbmsuamVgasFwcTiLCM4fLtJOAlmdtqlZESDWtpoa9zgqMc+4PNDpFHHEkXwM/1Na
g7y83afFQYqAPiutpfgRrygmKljexvZv2Vv1WZ/mSku+lYo24HfH5qXoIo/HBat/Jmz2mROZOqVM
7yzlrmNlbyf+I9l0bCyyr58z6wvj6tAHnJnHk6kJ4Jqnw1TZMmbQHsyYYl+1/pIVkdF/kIwlVojw
HP+2h4YjoEEwefzfmSNN98pB6x/pfimufwDcyiCQcBUVyELZAYyFwrVrDvxZBnBac395DZUV3em8
PjhZZk2+ImTPmmAB5d+U9V+VSWNh9hAYCsrbVf+d9p0iiyPaLDrw2nUMMmaTn2VwSM0kYk0Zerjw
JwfJaU/XpZUAqk7v1tLB8ovGOckbygQ1yweWohfuzZuo0Zsot3cc4Osvs/lsGT32iBlo7buFGp/X
oscQXfUTvipxwufa5DeArDyDx1MuSgChf4KI+mTOWaldqoP/KOej5zpD1jNUv0eyB5G+6W0WrgD5
6MMTKDF4GdQSyG/NS2D+Iu5/vjeTw8CpWMUZrE5w5pdmfAMs2dfd6KGPE5Ggv15Jd0VPunk+QeXm
aXewl9EibRs7iySfKfLcI4m9VY7c1R/bkCoY96zO2ceXVob/SE1snzfbov+Ok77nx7jkBVKgBZn4
Waj807L+p8RMWzXYSrhmr90O4PKfOujZ7PgVlpygjKlRsrmX1dkeplY0K6tNqlSDphXMC7UsVlIq
CqlaUpWL1NE7/1Ti7MwyzJuhYGMZQE6IYo54aixVECsv58Ih8xhSJny2T6zhk468lSFPXqFJFMPi
R5WlEc6F81m7fkBL4XsQul/2S20JH3sXjp/KyWehkvQuHtPQH90RTP887sqA+TiazyiqnV+5GR0h
Q4L+hutzOYveUCX9zXEbdMlLeeayTUs2c2qhN3xRMU48B1+MW7koy2SUhmx+AYTsveDjcbAd7jHW
NLgXFQ919IJRLQ9ikn0/lxhaH+UyfLX8UvDKGDuxQMPUSsfTZ6Ke0P3Cy1vmdRcGlEw9mOsUe/+J
ZzElZZzWoU8hGl+y04fomWAYwo8pTd0n1O8dJCZJyyngTNhhUHW0jxTM891LL7VIVUPSI2cyOvEV
p1br1trVuJCBPqVjqDG9pe09dCXpTXcUS8e5r2+mF9nvtoCoFOGg5aoMcAJ6Kn65o+MCrfFX1sWq
u+hXGp+yfK5R2mUUneqEEG3ON8OY5qo/c5bJY3O7T/qItqnCl4bo7u+oqk2EsgPYxAV/NgRyOHff
IArndpyzX56OFh4350lWiinF9P3QGFm1ccgww1h8EKK4VrgnKtsS+WMy9c/Dw3rKSXHHt6bHZqly
zlzOMGR6efDTBSNp0yggxD8F7oWGNdiQsy3txj8HRXDG/jvZ7+mIFZxVD+Qr9Yog1gMvzIfCMjF/
RUOMjtuVpx54vhOK+sjwEYoBxk1NO3JyIwye+BNupFoRMxvLigszSmN/CJDcYEKgYoDieY4Ynt2E
esKX/4CE5E3vNmYLVj4VYXGBfG/VysEes4HQtvP0Mbpj2HRl5JnRM3VipvPlK0BUnjRVR676zTNP
w+Q9lv6HbKwUcFHNyeQKqc1iZwUqYr6TJ/eaxbGt+SXvGyt60s5/01N8UeWzaNqsjG1xT4xWbO9K
hb6H5PBdmVNni3D7rX/rloK1BmEzZiCunRls7sbdklA3Vuu7kRrziHLuZoW4wexnogt+BdOz6YqF
4uBIomJS/LJaH1EV0bOcIzNM2y+iyxOJBCEasIfAR3a51RDTU92RM7fUYBaBp0ZPICclee1+hSSx
Pf/5HZ9dlf5v9tQhLWaaBuZk9eE18E8hBmpaVAKFOlRlVsIHG+JKh/djiG2yAN8quvi+gxGFro+T
u1ZZGt2pYbumX8SqVDwWStpumaJBnKycXBXMcZwarIAalW1ysnDAD69fUW6rekMQGxANsJ0qmze4
yzpbv++s//VyRHiManW5PFTKVToa2mII1/Z2b2RGrGETm434OCQjevDIqMoaV9Pd8wdksPfF2fvP
EZ8c1jKYcvLm2eFicaxgD6hP2t3jZXSjBc31KH9nf7J1GnRN5bc3RMveS46m2jeycREw6KP+hw2w
2/sANFhOfuO/zkvycQuqKOUtXxMGLgT7G2gP/iKtOHlcvVBEJdOkfGhNie72DyQ2Pv6+iwQjwH6C
iySUg1RLpUA/mWSFFTCO6xRfjnl8s+u5uea1wAtcSIaqWb0ZmJ5yoskjEXem1CWRkO/XXEMyopcd
8+QvK1GRfN/C6hOySwffJW6WH7G4KFe1kazTmbLTvccCwlIu9C4gOkiD61m/E95ugGxLN0PQsLJb
qXc0w8Iq+g+Q3NMl7OEfuLK3kYsFEIN9GNvoyF9ckAMwEQHLBQ3U/nZXJyZSjtaUJkDPJAh4pwwH
QLPOUtkzLL1pxw7y6mCl+v0dphDgC3J+u2OW51ziSqWo3IefYDZOKTLWquK01p1JWu319epnpwKS
M5aQyrJRLMpD+WKY3MFCPMLFWE5bCnVpY29yIotU1b830OItXcPpzM77RGFnPHJYq5lKRYJJNbux
t/vwUFlYOE6sputoHLrynwHm5l0FvNkVqqtSvng1LgvSukrG9CP0YN2zdnGSSOltYJKlHpHo4VWo
DBZEKwjWvFIJXTB2/GJcDag5CKp2cVFBYaHdXu3jWWKU95/qe+xC7JS6Un9ILBb+6H2Sj3VYSp8Q
BA3uTzDfgMQMdZlgy+3i5oyVkY86BNPaVd/ysZrfSHqSaZ1iSK2DNLH4Q1J+kJ8f2JSmZ3gJqg0h
HZt5zWL04p44IL0bVQRXn7wLF+j6Wn8sY8YCtl5/9h72lD35XOX289MNOuL22OSiRHb31WGpEPiZ
0QSNUjpX6pyaSYQnQS/Ua0Yi6mljW++07iokk2bucUZFp3FadwSMUcioRb7R6VtdnBPDTo6ncbWs
Yksx1XJMqjui3ayxgYxq8TIRDhni6YLHdUuT34gcVejgYN/KyU8uQKFFiSjxcEPMZFI2ygXp8LA4
prbmNRD/nsm0P/CpvBaMY/bpAf3JGDEG4H6Zez5F+abdjlPy6o8EdvFqw7S9dux7FaYm52MsTxP3
0t/VD3wd5che7smO9SpHmDQ+vD+1i05nTJGfLnkCcK4w2P/GcLL5aeIGUcdqYTfPRP7SG1bmmU2U
qr0wYsR2U8HOalpoVP+4LcJZKz+9/y5Q8HSqmxbNzD6IQDX8CRBYDlzmp18esX8Y3ED3OAolldY8
JPrhDev2PrXOodFU/Jc4DQMstRJsT0Stj5qMW3ajAigyBh4z+mtxbdQqMu98reFMITOp+RP2lhZz
SkcKFQghH9oxOehU6+O0ibZhzzwXqrYnIiDNLVg9FmoHakK0z7aOsHn3Gk+bEIaaEDMGnZGVBWin
FVHT8+t/H/ukl22JhDzhjoh2P+1WEqak7LYjRkDJHYKPUtDP+mdYMJgZLcQOZWUZKeH2/RMJVvqi
j/UzRo4OUI7PZgW/zHO/lggvWIcVmyqhzcOcHMzzEqLzSJxldVyfvSynmqmPEIBqhCzJZzQ8fy1c
C7cR3nSi8MBurzzkombHgK4wEOUGMG94jFBexEwxXHUwINT/dsVgzWYPccLh61Ridz66Fw0sn6Yy
en0tqKQCB8l0KjXgdha3KQmW07GEvBG5UINcd8cnmMhX/x/uKAdU2phLCsj1C6DBrg9Y5ddLaxGS
KbUtCi/GRwMoqTIiSnTW+ss2TMPM3N5C2CI97hHg/RkgojQIg6uRMVsHUhoqp98Wk9HjzDcFYBcO
l6n8Ty2bx+TkO349Fm7+MYXRfAJCAjopjdH3iiQiOqsB4l/A7IaXVENqBIrPC5zSyE7EUeJZqkg3
otDnVAUTdc/cKG5RDn1p6zz/sY0BJ86WccIjSP69pdV6HTcy5wBaZFCBbsv4zVHBhPx9/9Eiu1RR
YZRWUcB0oopmkIxDZJVDTt3ryx5Hk48R6H1hWaYCkSpAT2afpBalLnQkoGzOJ4b3cHj5bFY8vazZ
WJC0jH314pMxEGE+x0pzQA29J0s2vyfXmdbOIawcYtGqW9zV+JNldpj78Otwa0jPyd5O4b1dqz+Z
P4J6wt67d398jxLqpsgFFBz+D5UBovz8/UBVKZmG+JuoaP3wI1Jt7F8+OZ1B9hT1boSnXzl3p42j
LPisxc2+bfxXoNyRnK/3Un2PQyJobNdtn24zR60TYhh123JfrsyrP5fI7MSMG4oTdldlIwu1NSRA
H+7NGYvdwpOeVpuYXFehFNWf/kvBjOpbquNVPmzZSE+IXOvYbM3tBoiaHa+4pIo7Wn6DkwgGJjbd
Ptz8AOSfVcBQpcs93Rqyb00BLn2YNWJ5k1v+Bw7W+alsAA5FSTZHLT27kT27TcOzg66wqA25+5lz
HijPwjTa5iriW8UMajCij62jt0d3qcaegKkubxft1m3BdTAaYjYlKFelnwPcKcCjTPyiuPrkwQan
0UoyCI050JkOdbOIIXolPWkFS3AYGWupHgHYqjafA80952kr6RP05iRWIh2phVMaY+LP4Et6UFiR
gU1W3dAupaziuFtigrdBydRl8agjaMP7erJ7s1xV0e4k/LNGNnwmuuF+uaMS4uoYjqQi62aSHvB4
Qe0Exx+rToC/hKFDAUtetomP1DM3Zzzb4tXHkKoAaKTGmiSEM8Gu60rsutqJDAKwhexNBRQz8dNn
sQyKV8RM/HnYBSCayWR7ih/sKexTFZru1Zy+OQD0TJf5+46uAqVY0RhLKhiTgQh7j/SZpJZITDrE
UEUlgo2ZdhbczwnjHM7gm2gaW/L81zwuylR1+VH1Zd+70pK53Bbdb+j2WxgdlvpGOWtzuWruvsd2
ViZdlKK/ywMxZynB3D0HPyBHX9NKHKQRKwpVDlkiIwxwj1wB8VjOZITjS8EQ3KIOo0zC7AIhvL6Y
sABguOVriKgQ87jIKhONuKRvCJmasteH1a0hDQEbsaT8pHAB0eOaNokY3Ps0Cu6R6k6wDLIRvCvv
5W9yrNF16eFWbTxxFWiy4VMRBnl/LH+vp/bNhwVBTs1yn5wisv9UrW+dSYJJBUk75x7tTWyFiyW0
S81rchnSDFd9duXXLpmwBBCogFzAuMuUf4S0Zen0DBWPyXhY/tS5euV+oOC0ttwxBsNzF67m3g0T
ifXsX/nsLGJC3MlcgJ/qJ12iD6R/DjKNC84fjE+qYDxSqGBic3kREd0xiRe9wa1lmH4YmUpNLH/B
wtwjVvvaUCKngh69lMjDZhg6iJYXR6KGROnAi8qn/GRuJDclT4sbkgoBQ2urrW68A8hEfGrvapql
ajBaLAzyrV8dW/SzW4zsx8tFv8GthS4tyf6sTZlq9QduUXuclxZQ35fk1zRdOtkZoDfRJWRaoJ4R
Z5x8mz52wK0d14ruDTU3t1ZKgk0T9dFXX2PbgiqUFYkbDV8oaMtPObkZaT4B+dSUzFN46mwhd0Yd
mZVDSeKtd4m9k+dD5VYC25oexLLrDnEvTJAQXYjJ10IAnxxJ/QR1XjTQ+wN+t5+y37qxbdk2YEcb
1XQgxRjCcDJii5YUyRg/zGwDRkuKam/Fjf7KP1anypIWgE1fsmOpMlvGFVMLm/0aQ0qUGmMK3fSK
1ghWVNcDEf8cknY3ESFSROMUO2Ez9LxtBzmyDW4BWBlajPnX1X6CKqZKxUzNe03oM0TnTBrA53hn
BhAwkiSOafNSNhGzP3JHO+CefwWI5UaKKGJ6RXqaM1/Ibfd53ZSHgB3PfYN1vg0hGXoG3DNaD2se
kbytJITANBCxTKSpe45/XB7oJu9glqa06ntzsnXwSqtWkReuyaLNE2d2QMxBWwNxCrD/pA8vhywQ
sqllxIF90XAF+XNiSYSYKwLdmYaCTrmr7Y/Am68s691oH6NebI55TFJdKrEaPLhCqqOWGSs3/m7D
6TPg6tynNq7x70rkEO3YpDwI1j4mR1v0OGq77/v/g4fGtUAxZEY2gQTCBmQ6irmRXG/clzpxY49F
H89esykZh/70BEZN06yEVGUVVr0qAoQrsbvc7ycTWBY5bEpP4ZNCP/kP26gLx9Yn6enoivt0celp
YD2mwwXe0Gj43Bf4THpkE23ht/6r2umU11ZLwLOiGmaWFxEJWht30kHX2SXS9PIrUWj2kObDleH7
6PzRjJVVA2Xg/EUJQSVjcRAMcYSGT26JDlsb1dVH2zCqRI4RqjGBst8OEYOc35dkW5PWAGurI2tk
857TtmImCR2nB0RTweT9S3JZSoFWea7/u4AsDWQ6p9O5O/d7dW6+p/JYWQqGi4cAEOr1MQDVclH9
N8KKx3Ox1ZIS72V55tLXj8QGAKLlk4yCqjMjG4QKqonEhGNuwBAW2EMW+ghQadrvhBUnPqTQ+FR8
7VQoOGTcwXnuR5XrGWPacQGUnXFsWeBj9PMLmsyjUdgN+gDFvDm1h0ZkRPaGJ7bmQXi5Gz/X0j7f
M4SHdb/SR+//ktBWMWrr9xC9j3Al3r1brCVXhuUG4IlQyZROx9hphD3vMN2CXdlyr0o2ZtBLgCAu
qpn+bHagFaK2KJoXcm9pkJveeTQPgxXa9ASpRplgpPG8yaHWVeyjv5PVrBZIN+UDrr+NUennbiWk
RpwapY2SdYyM9+WdmYZNOwXofziGYS/Ksc+KpFby/bagu/5KixSqAE1r4XuhOVrP8L7C3W/V3SJv
ljDjy/r+xb7vasyAMrwgC9qO9MP1qtE1q1WvKX5eGxt2X0ZXMfXhAhB3/XP9OSEmSopyN7zLTmVl
6BCb2+6KXwmFZ4WLTDClFHclV1XlcqpSjmdEpBhYzhfllaskKl+YeGY+48oqh2Yx2IG8AKi9KfUs
aufNL2twhFhkCc+8U6hSj7u5QpFEI6/j81oeWUv74J6A8stEQvfi5TJHUFhIhtpXFi3vrSSgcJFm
vlVELVP6Zd2UJRkzk0W4B+46oKWd00liNVyttcGD64JUcLtx6U0E7ARcXYbvXvF9jz09pW7ITy4x
KwwaPfzP2JPYKWAJhI+JanISpLwf0v0nFHG86KEKVlIwjPphVg8jvIkJnZIrtx9xYFGgkiRpJmuM
VYpV2rApsz6jrjUqVm6GPh6jDQn/mqKIGL953Ymbe/AVB+8xRDlkikrOY/aWJwZ6qciXsslQudQw
K17zLdXJBkXk1/nGZZwQ/vIwvh2VnRBErzzxsDrOJy/V5UT7riIXlg5s0ofyBUOhHq8rEXslDe4p
kY4QGTJTXP61QhlkTjA8RG7ZiZWZzfd2DnqJpLHMsEmxOpJFAT1CXKnjHCl3HwD3kYC5D2Ho2+G9
WgZ9FqNCYAJZvxk2OCaYMscaAlFI8Z65qcVsz+hUk23Z+1s7XZqfUvh86Ys3cgxlApFEE96HezsE
Hbn+DeH7YyMXisDo8cP+lFLNM6oPPw7Wd015YvCICUtsL9Rs8rK7OKGU/ForhRBOEHOix5bGtMV3
f+AynRF1Xs52SuKQoWBhfrk6oR7ab+VqUbjmtsY3c8CPJt8npFE+QerLAW52TCFdSUrtUkOR3fM5
zi2vuUCUUvRIqHUta2fdpzrqtn3CRAtCFrjcZ/Jkb1JNepivRbmQrUKMX7NDukMGf2sohE8RO3DI
vsHpWa549qlfpR1N+0T2Aapy9CYKDqOZozHCMRISIDUzHm+3ZOM5dFoe2L0TcPkq10up0c3LTYV2
WEen45ZOA6Loy3a14a1CEffnOjnX/UWoe7plTOV+UC09WrQaTd+JsfG1CqTPJbkFDdz7jwwXvmNz
VvQQSwNB0LM7edlXJK6oeZXxs48LqWL3fK3eNrLgtuyh0yagKOp1f9A7+TcErY/qMbqCVT18HNAT
YmLqcRa9iso6IwKNUBbS3qcrt5RTb274HDEFLRYKkqxR/3BY+ZH/roTr8+vXNQ9P66Bql7d28B/l
a+C6yPK8wdTwNTUhLf90mlRkl3/KJyIAtSIXVQsL3cUOkVQKDcB9Y4sAPwosb6I5ov8m/0J0UhEH
/RBbOdgZtbg/SweRdj5NGwULNLjOuuMmEiHeb3B/Yw1aSJnY6Hu3DIcfq4OV/ZVBVUw6PCG+MzON
xtYh1111gPGBMdqUaFarCM8g5Jwhn5P35T5S2fHVDKOimqXW/emcHe9Oe/eVKR4j9RHX7k6AvmDf
Oybn8Ui0v/0bygzPW+PatS5sG3rI0sG6ZdIvMI7JLD9YdTX+yD17PMMqP3u7/MTGNxNmEkGv8Sdk
KC1Ii5V0z9gTi8hGKGVo9oWBtRAdVygpSlGCYjOWbsvtKI9mf/wK5gPooeyb8+fBKgI2wImwbabz
AxyWezYX4YtLum8gQMro2G+FIlF1JQ/cl7p/MqWyYYeQOO5qz7RYDxb1f4cgg/dHqgYdBiJyi7gz
NJMeC3DCzm8ntaA8gX3OaQMb8FT/YiRTVSn/2OIKFBfeJAmPm+yfa0ZLjJ4REskpqtSY/01LTk6g
LDL63DckPy0Ba/Gn7szHVzyfUXglQKFEI8CcRImkcS9Fr7+jlnGQS86FE3SVmM6v48AioJsOJJxs
TMZSeMbbvJCNUJcEpfjprFgKCWTQqWFfZUBoJAyUvBj4ZPwO9r/Cxd8kqISpP6fFi3trDiU7H+NN
N0PoCxvotA4yQh1kfqnHtQObpoPFQ3SdIfEgsgwD9E5+K8oopbsPs9mV5Rs0ENkicShWLy1iW4P7
2lvOwkqP+fWzERGyRP1T0c6a78wcDxFP4zdxbMbQBvT0A3IrR0ToZqd70Xy28SbasFShyt/3+/my
xjdekEIG7EvPpE/doNvgvIUeuoYpaxKIi8NXL4eOMUXXm6As5AYG89RCHd9mqwWQPmVLqgeCS8YV
mkalcurhZZUCHFTGpYd6yjh6BAQlX3RTlsC3xYMfkLwhUfr/EtHsNYZ4TvM/NdwYDPhyHoF61yaf
mDHa/e822O7HLaYmqmGX9qg4ew4JZOV7kDSw3LsYx71P1lEkFuolUKeRGRe85AGLenf6dfj39BrO
yElJzLqsYIG9EdJsutHoJmUVOgW6gqeGagqhDiaH1CVEnojtpZ0FN+yHR0GVzS41pDTUQJy7a3WJ
nQKaYyMoJCI4WAifE4FjJp6gRypc+SoyPKoUT1Rn2lmL6TMsMtVUbvlsdRyNtnP4JhCxf1UKC8k0
K/OdKEKSeqqWY9aYD1b3r9VpCOxeNJ3ltvXIS32F9PFpj2VlIC94C4R7HqX8tq83SxrmTP+GhBr5
Ev5FI5FRX5qXPnPMDBy2KUq9O8LQrBEY4a/v6aJftd34vew3Dqyq6wargqYD/aTykcV1s1Hq9/MU
C2iDo4QzCAjEOCgwTRAbGpRQ+8iS2un6m1oeo/B5zKT9eos6sz6JMpKwwTwFP+F8g0j8GNzXgED0
YOTnp+7lk+DdsQnskNtF0XAMklCTquhOWpa1/Yo7vOqnDBie8gt30m6mEYUTw+hfyc2NccXLujcl
OETi1qra5fbbugQ4QYKy0WLQ6N2VAUShynxx73RZxnwhSVwVAeCn94sraF3kLEqtTx+BbfR1Ch8t
9DJaKU/K9jajxwCTSdt93rykMJvpdo6TvgYHcUZ5mItOY6RPvjX/KPq4tEGtzs13McmzMr0zPmno
yxaHOeif3JGhhu0n4CZKDqo3M9sWITrSHSCp19iuE8JgM292AFajVD4IY24TDNCmbxi2tga+IfaB
yFdnscYiWa3Tp9gAIqc/m8dJ9L2pi+H1U/XyDfNCuLPJ/51cFv+oNJ60aWHlWVd+Rs+qZEoF9zKz
NogGAFTZcKBPiONtfLGp1MzdbrRBbwLJZE7OdppSZAR3448QhW/5Tm72PONu9FOoNoFJdi5GmWjS
oWCpXCS1dKclFYOwJ4XYUvnPb9P/MpwPG2DXSZaKNrET0rdKbD1wY8kQSS0HWx5bnoqDU9jDIgrD
xtkFQROKq29Uk9JyeOk0J+C9MKQfLi1rLuTl2RvKNS0wrLqd5afgIczOhR1PbQpEiwB3vADOkjm4
2aAZMU1aCM2NCRRbB7+Oe9DMusabfk41MnP90O4JQRY3JwiiMg2KC1tcOxbyjM5+ANXkfPk+od8o
KmYYYR9cnznpQQG+rPCpYqJWUEEqm7bkGOhsSAL9BrPXofq1x4NdTVyBAOejEd/hbLp73zYT9Ejr
9iDA/R85noavVP+lGUEV4e7ukp5V5fxdbdf/pTFL3Q4tkVjalI7ew3C07I0bpuIqbQklN6qG1/42
/oya5nlTq2DXgQpCsYid1yWBjfGlVU3LgL8r40uxOGTgqKbF4PVSUacZrl03F/9V0TqZEKJRnvZ0
nTPKM0kwsk2iOJkWtLfigUtcBks+SbuOixkzNkvBnA8G7wa275dTV0Nja/MLbl2dW0rR95Z4Wiui
gMcZOUFPx1SE+yxmkaaEkcd0+E6wFu/+7TXz3LpSiX9otrDCPH1w2/uueaJE2O/soijFVquyP/bB
hQOpLDMvy026aWaMLG12114CWttuea28ECtw4KrDteHQyFqovefuaQKrmANhAn+HiBPP8JqGbKN3
4pKu19rs1xppkCwehZp12TofI8fyLtWXFmQDYq0IZJrobvrYOGggOq8GZgpxBITCjB0avjl/JFgP
a0ViHy0e5lOQkNvcqszCQSqYr5EtNRcHaMySSikrBgFEEKMJnATjdwpv1gqnSiJl8tw6JT2pfAwK
b9Ui4B16G/UxTUQrsgbAicNCd+/YEKUQAq3A67KBJ20Eg9DqU13DxlG0U9E8bE9qnre6YpysCqV+
AZBpeARcyOzJrte0LzT+9CVPv1v0xZsHj5sCuX7SMB1TihtwYdldlYjL+Egitn9X1YIm+fgb/wGC
QL0srFtcBJwUtUhKmUhJ4NnT57NiR1hq+JPQMDGpoe4aqHh6VfCLiSohsZyfRGVI54fu2HPdypSk
sxM7EGJ6a5jh3XFJZyRgY5yn51vCwhq5HoUAAEUKoqFmXYmOwr1tp9wCtX4UVfRvLoPEoyvA1PAw
I+dyshbJlE01zum4qW0VolwXfQdW8XOHBjnrR4z6q0hz/DJSf6aU6CyDg1f3OwNvh2Lk+mn7Iq2q
RjGnXBbAAsCwDkF0KtRUmq4k8PGzgZrazGeh5RD5Z27Pt184e5Q7/GDW5xZiHjdMmeXQrjdDe3Q4
aeMN91paMJzfryN3ifY9KHyO4FilTZVOVG+drwJ5/lk/kGj7GwB9SWUFxLsDhQTKYx57G7CawUYZ
METU8EzmYxW3FP4dqGayMgi39O8P3nDWl86eYwpdYgOLK6g0X38rUAXn4G/akXQwbXhl2HOgxbTl
A/hwwbpo16mA957lFMwEp4YbZglMUspM4COEcZB51IT3YPNtKW50bH8HDPSh3sCmNPO4OX9a8a8n
/Sx7OmAqa5p9Ob2pEFF/xqAgAjMz7rLpiaY7cFE4ZCJ0mXT8i9SDm8noc2tu0AexlJeDZOJ7dQp+
R4HHalLu1lAehNI1C8ecZ2F5UrZPWH/OQTXjqRDm5O4p9ZmgJmolDCsE2+6Kk5wp/6bgzO2NxVEM
n0LgdvAf9m2J8BJG3kG33So/UKwVwtPA3gwq8jWeTMEPmhqywXe0k+6gy/y9NkUKXIPUJgrNBknV
leGCvWbQAZaAsSxmH6EHI7Bc3hze5H5C6JQFGu8RpPzJyLkzwaCLvMt9dFQzYVQBLXmnMN/F9hQF
tNxiuV6qORjxdo/vM3jq/gDucYdFk+2zLTXTAvBuFMo/04emK+J3jbJg35fdUMjbXq5vtTEPQFtA
xJ02bLoLz2zdBsUjFE2E1MbMoFqoW1O0lB8kPUke17q4OUtO5OxlEgOsw4gEj8bFgCDu7iiFsrI6
7bvN2OPs9PEHwZizbd1m3TvsjPf6HjlcxMUwXK10ZwK7xGEeAP0flZsml4WUq4cv2lWhPG8wgo7N
ZGeiTuCOS8UMNV/O/cdZZWQlyna89jCwCb+pTYmnYmQIhb3Bg5AjhTpoYOAG9qdGM8930nfWDfJ7
RH5Pv6vgGqA9E1LNtJOfiyL+ezwUMuWF4WqSVFgQA61bAK/VTfBEwFYrtfkdzJDjC2GRBEcYOE3x
peDAqkqHPdqN/mCcWmAWfCQatF3iVAfS/2tzcIjIwnqt2rpeAafPwSwwV/jDnMUGirhNhJHWFdMW
TgCXNtdy0HBAq8xEk3c34TbS4t2BOyEVMs5D4WhnLJoBMNiGMercJcg5Tqto9y70KBCgE4bNkR6k
G8F4xuRRKAkDijh6h39oaCbPrBNCiIJFObCVAdf/XpYfLrnp3kP6HEe5XqO6yj4EA8FSmQr3u/CK
/3jWCjd31BfgTAiByWl8A6JsEsgZUPkMX0QN//0EZ+Vbe7gSqi/zpvMie1/aOmdf+8eI0vJrzfY8
YFE1FiZxDZv6kXrA5szsg0ey5UagEKgOVrA5HdHffNTuJEuH8cv+Q3FbJaKW0+McSzrKlQ7hlUfr
rv9Tkg+D4eNHWZdXeQCYIQ1PWJ6dWmhhx2S5v/oAEeXks1ZOiaNfEiCV+YkcDvMEYCcp7EeJAeYS
bKElbVr6iV6toTXovmX9bDh2G9fn9wwaUsKKFqH0hXWT58zhQGnSn9ynytroQhSOqsLhJhvRy4As
Pw662waWGPOyRAfkjkEZXbraMy89h/KxJko0V6+TRn5pHAa58h9hthq+VhPuN5HnKwOH0d3UXrj8
TcmXvDlpO6qzLUpweopdyh88m1CeQ+xK616wowITrGj7VpOFylS1+xFgzY4iJQpIDp1TTP+slCop
5kErl0B3t0CH+/2qMRy0LIT+WZg0DRfZOLLyO++54jVmOfinzRi4g5VD2A7fU/9WBvsm0KiaCDEE
W7oHFgSmCGX14b4C4jmWHliBxott+qGTXUSq1AG/DdXjMPvKpnKq4ylGfFeIwusimyd45k/LW+nq
y9rZyQoojfjjcJ4gINoLl20LIgzDwzhpt2my8uAIpvV0XKA7RqEfglCR76D3SKhcs1KQabSzhXCt
sy5LCrr2spk7fn8cZg07+/s2OR7aNgfNmkX7VPmO1gSREl6Gu8qpz4sVEgoK8PSW+FsYUh5OWYYn
ZShWof/njIxcVx4sR7etv2wOPM99OVxY4eo9AaJMVydZrOhBlljRoRztntYYXEOgwpj4790DUL9+
Ujjru5j0f+nVReAqzPcAUS3BLRNAD/uoUdgv4UpoDuxi+zg0hDmn3iaUUBOOwxJE51Duhjd6aZ2c
Qw+h45rpTb4liOqHii/KJuDkcDj98/ynp4Z8XSOl3JRRd1VOz0ivb+4U4OzBUr7/+luW3gAtCg00
MoVkvz/bhrSO1yjrWif3gK4868h+QrDrHr6RSGbftVzQaRWXcWlzJKm6ZKgCn7N0FG10GkEkmrXR
ChCJ+JplI60dhRFB7K2W5Z/6SMnTzmw0iXGPTiwEWGc0DPfH6RGxslVhweKZDRQUyc+Oz4CCMKzz
XUPlbxQZoShSu5Uj7Fzpa4kqaK2072kyX+jufjEu5MKywk8aEHAqp0EWk2O83ezQMPjGDwl1ejJM
SCzBiE36eGi5ND+gY596XdPN1THESHWVDOLZJcrJHZn6jB5H0IlM9rqm0z69iCv1VWXRHkeW+s3l
kY//WvB9brbVCr9JE2zOYIlgre5OKDyLhXIHjJdaHhNfBLfOwFOgSFEZrUkBbbhaIvvAV2Ah1L/u
C08GlQXF/aip0LYrjHcwebAkkpxT4gvI/p7b71+0KsZadHRU3vDWZNrNmkxE/sXYMy+euPeeVCIg
dvOn2rBIwyaNJfouj0sEgvwWZ0FUzBapftp6S+Ar7+3cijPIwbnrRQ5XJbLv1WOccCD1n4nEdNG4
3+CxL9teJKOoawfJtOjIGMzHDIyw2K2tQT8+tQag5EQmyxQFzTSMg76HwmoIQZIoWQ4QPfLFg8BE
4Um/25Y4UKr3kqn2MM5iFWNR8Q/lbuU/VedfJDnYXb1LljFfSgmxwlRVdj8o9T9UtccQg3won/4L
N+w30Vflypb6noUJsF6mV8uPKKa6H2cJTjU27GUb7fINpCtq66GkbySyIccq234wL4wXQKLg74/L
s0ql59Nzifa2bxsWXTzIOgfAYM3OswHqNKuMv1qCjaDtnhkLtsCqOmLuxXydrozp7KkaSow3Au+E
ENWxW9Gyqph3lJ6HFz8jP/l0z8klPvwlKpqXGiuJ2Y/ZnlJcurYB3Kyr4bYdSwlOakj/mmwtXDcs
7XzHrFpgZMUugL4aM6qbfT6YRfAcT2jhf92LYxbly8TiQWzFSpcdCzcNv7+ECM3B9SA4lI/GAP92
bLC34I/1fP7xyzWymczaWkQVUGq8DW8M42D4FjriHaspnClAIO/9/qT16wdWtAahPJFhIM4XidWI
TTzbj4XminI7QcLL6TGkUvAivHFuoOT0qPYhOcB7jFondDt35kWUznjwHQs4frq6VwjiTTHRZ5Fy
/YRQiitnBfaoLcS70VGcuxMghnOLJyziBnSxkZVckQXhbGmU2wWxYBDhZPfQUwfDzWjfeAC5i+0k
rmJC4tbpNlHvA1cfr8symKVFAiWx+Qrh8QHMFkDp35j5yNvG73yGWtFkdX4cR+xvtECFam0O2IAU
qMhd/odwWp2aIGqWylG4nqLjk/fjvcXETPsE0+GYLXLoawtgKwhqOQCCj3uaS5bBUJYKyIufb872
f1BxYRK1iTTy9iaZ3NiEdS6vqPPHEYZntPIp1wB8QMkFPU38QomWTYCNFOZYq4RpX0fDOwLoB1S2
pCKd3b8NhEhS9q0I9XtKpgx1SNFPb4zD8WIzrYwD+VOrGzu+RZzXicvfsIkbWz0J8GlJXf5HXVb/
wkjRoFTnKb1MhSdgBKrcZer1+D5iGJcgMVjRyjMIUuqQC4YLz+4Bzk+cwyH0MEso20zjAMVLiaGQ
dWDY+sLJCyFnuVMA30gi9vkQBaCIsmIUp/hz5V/jI+1ODi6uaocBNnwzcjYrUXbiipaI/4/neSJK
1jEWn9eRSYg1tAYpN3UROXDhGQ0jG/FleYaj5mOOns7CVzWkVd/M661PXADMZmTKq2jtWGQDvBYv
3B8KDih3/nI/NKgjlgnfCfumAYZ18EfQvNCvvz/+tpOaMnul5ynx7N+cQ8rySEBWK/nklU+HStx9
c8hi6KVPm6izRy8IfXr7UN4XKMAqyBqkt3pLeU7LUZM8GYRIL8v42WvNerTLSBfl/yG0Kduo5k5W
pw0ReUb/qg+IghhamhPxI3w3liQPnQGlpCE3KZRfe6p4xvKbE915TRzz9myWByu7XnoCIJpPhClc
4OA5mF6Y6DkgVYzh5kj82fENZCkYwvZdI/mA4yIp/6wxvmoa3tu8wvX0jli2hMf9ycWgGGGO5Qij
K4mt2hlnkSfh3vG0fhbO963SeChAYrUYB5NaZ3yZMoxGS1dy8vMD8BL11IoaOJ8/2Yig6P9rBYnC
STw+LjNuA48m3QFy4wHk4FO7o8w3Q1L5ujNjWCIXKkNjh14uzD59kP+NftarLNelTR0PgoOqsoPe
ZWInbT8J/AxQikhQbx6o7Kbyu6+D1wIQ1M4463XBMq+A0tMRE1/LXgaAyQq12SPuz6+7MhQOU6YP
LG5LO/YD+XoHI8W43dVqKY0zga3TOIcmJ9MM3JVrKnD0Fz95vuMBYgpqeXuU2OoPv2S5Fd4rPPw7
1+3KjkQkXTqUV1PinOeALLu/iZK5haiBqHcU9zmMlkri1o6uWE1XNfQDmb8ruST/E5PQzXNrf4Ew
Bha8K3Ldi5f7zrJ+rPA01YzAZNNwFi12FsLtyY5FyartO6DOx9+fCHWOpqZoB1zzw9agzox7oPIM
LCGbTO8DMLT3DPE7K2DE+ofZOEDeqYhmdSfi6XX406Wai9NUduqGWZ6PZp9zv1AhQUJdZtLt/Hpo
jtOdFxEALpAv9M198KuLH4Zn6YdweSyF5yuO3yH4tbL2NoUBAxj0CuMpNeON/92WYZtmGw1SKsoF
3juxnx8TB+WaRHjHB7InOzEHVxhOoUbd9h/ti5vFlje0N/G+2VgfbqSk5COTHPVdBZ2/OGgRlRHK
suwMn/WSYSYZp/dRD62zD16DfHBlr3CzvH3WkQGvoe6gClE8fNjDRIXzb1Xb9WY7fgc31vbNg6y8
yty2GQLilkYJj57GQo44b0fB0IX7P6e6j3/APO08fmHrOMs8ms1K+XgMlgUgpHy6nPeC7Mg6gWSm
riJqkQJIQonKnWYdktxA6/94tQKiQGWjUCfZQX5bsrhlXiWFQicrDgub61cL3EecMBzCkxxgben3
1ub8YMV+C389inmKjXknNmj8YJNDsHIOOj792koar3PZsejggmKpBy3xt64Crw7WlGQnKdqFfkgq
/lHo4S3DkiPEJS3bHsr91z1exOyxawZa4vLw4AL8jrOcwvRRxxub+9QVEeywbVvxxAwksDDhHEar
aoPO9iZqgvMWYXXK4Cg+zOELIMKupcJ38wvO2VYE1A/RhGkcAJ7CrAOPYFUrUAFeOj09YlJja1wa
rPrtsi8JXtZvKIAp9UablkYOKxw7ysx3aZzZ/eW0pXOEVOvH5RRybVNX4SkTpoC2ze/4//HZtrb9
33v2JpPh4/H12/CrmPxzSiQ+oB+oOq2ITOl8ROVXQbyDms19I+kCuMa7SqBfq8pnj5oCu8igsajT
ENXya8Gz889alLh+jwbkZzYpVqMZmuHOdzQ8S62JQrFBKiF77olmjBOtnlT0shuBtut+ZA3Xe23m
DodZmlthTF3G/8CwLZk6uDs9RpK/tmM0YuQX6aNObEG7FOvqOpXPRw06yXjye5rs5DwqWZ++9gKq
G8PZQBPkmfvY84DV77VeyjSsXiLCD9Q2QmUQ3a/jgwfqy5AReF2+O3ZIWFqEtb0qzxP7it1lICCg
iaYRoj3mfOdSNOR02wqaSQ+WLmBIQLqx0oW+fZ/mPS8CFtYw60SJxPlNWbAebv5RMggomBgqegOn
aIstAWBNMFnbd7sKGKZuFtIKedSESCfUHelqnTqHofO/0U3tp9nV+i5J8T+nnKlYgSs1qnWhzXyh
FGIuwLXRc3OaUoZkfzjr6/N/GO+uRoIC+0Uf452Zem0RpvURbAgxs/bAf7AWSqQr/Q9cqtcSMEJw
PAWIFzwkRM7UiLoNIxu/jrHtZMkE/7sGANDbKmJQIwgpMkOTPUHJ0hiKTD5khMhwbtrlB+dnVCp+
AV37eBJUfbdZUU4/AwUTVMR7dFkIg+z57sUYyv//+F+O+q1jhNGoY4UZSjYDTOMhc6YsPAu1JdM0
yWjCGZPKcjnEq9gBTVtIyBnINMkHV0P3DY+HVo7zBV5Fcp08oBK1KrB2kJSDkwY9hUoXhK1gLc7o
wsiJybp3U6+8KiwsZouax85Id4HUj2P1pDytUr2cuhHNFQZwh1zH3d4HEN8j1t3KI+rpj6Dgger2
MDYP8bISB7duldUqkNfPz3Ir5G5ESe8CyrtP2KvUswcjIrs4TRGc2FdrNTErg1dqT/xU27ZLVhvB
uHCAoH6R28VcUgXiGK3HKOthQbBw9LSLm++UwX0SJEdlSScvUzr/H17TwVwkR3RVJJsnWkPebBph
8RH4hplHPEHjvOONFKdfs+e45uDsYP9rDNqxzO65pw1/Y0T37VOESKI8coRUzYpITwQyVsMqXgSu
VXlNWKuYcDyMiVaMdbAFFXxPOUZOfPFi4+19diUKbvQhMbakMRoKto14loZxQvLSbNjrGyHMCoBv
cE7UYI4N3F6xqEK6Gi0Rqt2tvT3Oo791d0U+1nQ3ARsvqJX9F2VmX/3xAmLLSt9dtrwLfa9XB9bo
6eDNHr3kBbSmqQXSlFzVcLU5MuQli8t1BS3qsnNC1oLIgjit33RWDaysRAvfRZPHmui4L8hyNaWn
jlzYmrkJ4R9MWZvwAlmTAsfA7luFs1GUKZffdcXNpmodTZaX7297Mi8GcWf5O0CrkSOuOsa3RxC6
+USv5VfR7gcwqR8X34nisVUmdmE17BFaRDHGwB30R4RrXtTISxqKz0QgOjE2H5Q4S4B00PLKUiGW
t92LwnzFmiwBAv8KTY/QLeHXtaycVqxC3mW6Xb5vcaSAnx9YtedGkBlD7Xm1IwaRpMpELeg1mjlV
DgByiP+0dwLlpDbNtxA8oLu/7LnnJ4RJwqXeftOJZ/dvND3RhxhASeOf9YjfRzCFvtsFfdTga4KF
cdz/uq+cTZDR4KxC5e3cxCyrExqsEve+/EaJJGMHkZHlA2p2sSH1ldd5FjmOs6xMKoxY4Ng/QLen
lEi7VoGnEZ8ZCwynC5DsvnPsgvA7XIvBwTCadnhnsNWR/YFVmwmJip3CrNlmGdqkvggK7CbN4S1M
xpP7/fVzYqozh/JpBSBXb8VE0niPvsUJmiLDMvwYcs1Q9sSA/JLTVG0lIZHguG7N3aDgoflryA51
bIJRGI98thH7/ES9vTQvLXO4tu3ymctKd/eFXZuYOb7ftn0WHw4SEac5ULXeJoGJLWWOJROlskr+
dgNjjAC6PwEMaUvR69Bj1sA3tdRxNViDrM9ko3/PXgvRI/DFNVkc+nNkgFPLBykyVJpXFvqXyOuY
ZVzdzUu9DPQwTvUj3KpUhCQVfNlp9MepO4RGDRHyimzyvWyVH+rmpCaz22qQqQ+kiLsaVR3D/ABR
9KwiwI+kXYtmbktcft+2u/k+GRpyN6KEYs2obv4wgp4W6pUF05uGq5QBPrCIiyziKhAkyXlKWeSj
6HK+nebcKYwfKFBPUvqfnn5d+FmtCuGGk+eTqWTQps2Ce7Rcs0KrXI3xtE0D9pXZpsuMmcU0SUnE
ueKJHzSA+bXgK8iCk0iqjsH2B+7THOSZI5RhD4ej8rWxmmVv/O6bBAyoTgPdrxixAI4daql6ZKLD
UD8+gbaF5FsxE2dk7mdkFLbzG8Pd1GrtZhpfdBblbohHMMkXGTjqkYiFe/tIvCrwCMli6+Mj0WsT
jYS2odhqnDnUSWhGjWmbRqE3KTecqSqRmkV54vUNcaANuQx6y+E8/+gBZRxQtZyGzqDuQZKfVIhi
OrHKZhNUWb/IuWdSuO3YWwaHbH+yODVeLvYcHVRY/Irre97IZQ18HoKdALn9RuDN7O6JB/t3VyxT
4tYFdkBptzcoKlcUfV2vvqcCxsmrsvYgQMDLIhLgUT2U4s7PQN5AlXInMoNn16xMbH9lZlHHzg9q
6pKTwwW/obCA88pYtlRrbul1aPi5DpQt9zT5UoK+D0gm5KmrtZRplxGJtrYM5q0rOx3BX2L3MtFg
1o3/0SuB5wcLd/YJ3sHKUnOa7dNfl/fz+S30kxqtRRreoubiGLLDIwT9lHqMnt2GVzEEBfVuq0vj
ZUr4AO+njVEmPdqc6708Qz4Ib9FYiz7f1RnfYWI3q/6n9P5GuzpsZhTttssBn1e+tzgeLS9gt8a6
IIgCa2jeNjLHgjPtdKap94B5suFZBgEi0d1YwqvNTqAhCjXff2YZUQ4FK9E8m3Z5+kRBNTa+aW7t
C4hVXuWm2UeeTR1MIsVzMu8z4cWMBzQAKmetci6xiDi3M2//rJ8CTK7x97vu8SolW2eZaaZXy/iX
MftzS8ISoxpoDeCrz+45C28Pc+HActkRgeZvNfNAtIQRusnWseASpfEo2shCpevOKdR91QNuJrKM
CB5kv0zvqCb6CfHIJ6SjNaP4qSLjST4zzRoqry6OeXGHW4u+jCw3wYkQhBEWMV4cQVUoKiW4SQZ9
NiDQ2nRrOrI874NO0e9wN1BP9NdG8xUoq6lUm6M3XaeKZ0lhgwLarz4Ym27KjsO2mZ4Depvy2Sox
Y9FHLCyvpKrzqfBBajj6X/M9pkLhziJiURoMJbMGuwvlzdj2zE3GDEH9ueURlvC43mNw9/xfpD4R
hrZVlQcUB78JVILICf/4Yw5zbuvp1f8RpNxzE7MTVINit9sCVniczLf+Jr6xzU6luae+luWp0B/q
WnYwnqKpgiti/CSD1ys6gK7YHmOaEehzPxj3brF6ee+vvq24IrVIGNM+oMuNLMg78qwu0C7tMdsd
t5215C/svhDZUVtAVRw0juJMtqTw/pERQytF781OTxfVco7msooe1pm7s1ZuQqPbo+7jue4jag2P
jlykjTr08bb+rRPblKJ912apPwK1cdwvyrjsUWVIPXvZRcgjvmw65g199zPtTpAQcNOFgj3mbIfp
BXFhN/Kyhouw6OUXTo9r5/5J6e1o4VML6VO5kkPepdm+1zQtkDceBZi7tXTMm2MwJvitvcAK7sx/
H/1zIfClFj+uq1cqShaEuXKDthR2L4vseVb24noCZ+bjtetvC/fv3FLOvl6pqVEEABiB5Vf3+51m
wappzMa4z9QBOdMYU1H9qwGe0TEyx8i+hNqUw0p9uGl4vq9Xsqg0+DioxLotbHFshbZFDiiITsRC
PGjM5M/3zy0tKvrOWPmQI497jhmjPhAh6HvlGQb3ude1lRhbC/9VaoSNY2y8IshUbJbx0MAZSLC2
z10MA+j7UdLnsd011Y2IbXCGTydJUNl8Z4rCjgVTceEqmxjRwmMNXuhSkp2VjZ4VTVFLXV4AQa+5
r2YtJwsFlNktKA7VglQcwcw+3zPsNdo9dhIJ5nz7niMmzyPGMGh8W9nnq7HyPQWMoCX8gKJsqk6v
yfL+U/p1kn1EiAvcSd/1z+VhJqzWqT+eBr4E4QjiW8xL8mdaaVeL7aUOg/eVqx15JZupZXLdV66u
Jfby02Q+tLPS/uEJMq40vi/Wm8FBFvoib8Wut0arsOimvb3V6To8J/LJee+m3koXHvoECQ9CBD9E
jagD8j6EwoTJGVzwrv77b5D7irgCTTnSlTrJ88aCIjZAyhJGs6O7nVGZChR/eFgP7b1RJEgup+K/
DRI7echrU/ZzWg/eCn/+88Zs2SnlvhMANWlhH8z228oRoRhTesRHnDBvzt4IhcHC4v8pBXYj3mFt
PguMdbVgwCim0TzUQD6FKfoopeZAj7hLCaohTbNB0Xh7KBjRCO+boDsBBnS0rsGplyiY9KQsTuAj
3fxBJd0vLxHztwd7mSjipNTfUjFwhvJiXmk2Xw9NMrzaPKBIXyPqg8wnfwVjTIjxHetXogINEFkX
MKjeaeN4vDhvwxMGCyaE3rZMeB4YOe2ZkUWyylS4Zbi091s6ukiy6xjkING63XRUNP8rJW41oxrQ
jDgSomOa0DKAThbcbS3xZOuPgL9ypTpkNcWNv2N3fNUvfBKJ47XA748PxnPBoI+prHl0tuKJFlTH
NNF1CLObDJ7yji+wiVwc7WJin5l2Y5n+rhbOqd/zOlzMRx1kgFOcyzM2HqIu/uG4ysgDPT75b+SA
0aIZPzJVpMxs6rAF+hs3h0SmPwFx1brJ8qfwUdMiSdsw3xeFHLuj0BNc71aEZzy6TEjD00BswWf9
wkCFiewCmmnB7WFIaKF3yGclcNmn1r5p98mYELtQeTNprpkBPlPOAbbOyTmPmC4EiJW2iTkZcAqO
np7f0/5rVa067VXHfSX5Fi01uq4sXE0hYdg21sZkfyBtBZ10HVwmyG9zqDPT9RphYytACjHjzqKX
tG55RW1wdhw+zurigjI8A9h+aTueRsdkczuX9Acj6ISacLlvFh4UDEPadXN3tDpnVfCPMs50CXLK
QI0emrYnhO6N14t4uM+ije7UYOPW4razuFdejvt3n3XTmkZU2+tKslu8anxks3EXub2a8Q+F9wD8
tV0k8+gf+xd8X8XlNhbb3+vCK/rbPHH3ghsDVte94piozqFnEwCyDPJWY/Dzsq7ZI9VsTDz+HBCn
Txssa7a6+94K+wYHYXVGnTz/vYvsSIBbA864lMcNze+oIFNHmlYdzuJPTro01iQxqTmZ0LI+wshg
0AQdvEyC6MdxATfTgjJpnRwiCZOMfoDlXxGD346zIUzrqsO5UkVtkV9Enow99Di4asDGaLQdN955
t0MCUKINl28qwqFh+ct/u31npNDpxUJ2Xom/Xu7jQSs5wa9A7ERSCOBKF1TgtWFofVf8pJ+WRnkT
YgRBtIKS6QRes5EMogBYZmljfC4FiZ9kFoI2mztjdp6Q1TJPJqyFCeV/hbglUPWaMcD2zdALjfhg
bQ64VqGKcwsMjVgzVdRRZ98UESv1AZvLvPDZkk2wYV+EWrndfYvim3vt4Q/VLK8G0B+aOUB59/9K
2nz6Vsq0Gy5GCyBMLoddglxxJYhAmkA4Le2LZIWXx9XQ2ahnu7BJc7oCZXyGHexvidG7UrMnW0DJ
Qp65FOjfZu7FPDNVDSI/Bun+SpWJLDKcg3t66Zn+DJXxNbhWUi14C8maiQtZQboTrPcBoV7wNJIF
f9c1nw7mTrb9Q0qzZFKXO5rYYmCUTcVYqSaexpXgGs8VpeBNwStyVuc+WEwRhUb8h4JRh3O3qa80
UnkxkIv5J2z3fiV2h80/mPrZHbjGfVZMEgVGIJtLKvbGEFLrvwfA2QeAfrrLtE2ni080z1TLVfrB
tE88H0FINQJwboLMkbl51laSMNQoJEqGYDx2MRa7d+dod1Db6wq584D6fBmZWBSqCzY/bqyy5QXI
DfyD/ZZmx1MZmw6ix4K2CFX89JYd5xL39eV+ZtuvXe71spNSLTsOstJZx5tb+WFkwyXft/H0Dxbn
SinqFyRO77vqzvkXGkMcESwpNwA3i/xsTl+1ZHdun/k6W3zBcRtSN7YkO6PfH6LDuvLGdg1YtCJ/
QEC1tMlFCu29MELfMxL/pIt+nHIXucW1VSe8n5Z3dUGBCQe9PvZVIl+w8vxtkbUL7Fsob++vqXZ4
1+vIFDjQcFFj5YXWlsfrlELDE3DNZGTjEWpw8b+adUnkPNY9KX+vi177wOuDLNEHvIKHfLe8FxPB
28ChuhmfACO3644r+4hhxWtzT6LRP8t/b5zwspozcA+r/1RWpj6CDedqnxZyp+BYQnGOEINqNHfL
Nv5xdv4fvAKeRHp1AKoYnx6tjiAKf0Xcs47iUlgaccqjTF2k8ey5nuJADJUUGWIPDk7WlB1NBQk3
MKO7tmIRNLIGuPnccbrWe+c2TVXE9wZeaRMkD94UpSs0Rr2ZEKH955OGkVsEVQyqDs3A+A8duo1T
jfoKYUJIzD0TyRwQOYsiPdfHmLLkGMNEdAKNJ7ka2xAUDQyZTHEWzglvz77H67vCrRNwDqp0QdOS
dq+R0UOjjFa3BoostSFp+7yz0+PE32CGmJBxkPJouOo/+wpuhx6lSiMx2Dw5+SOI73UaqH4Yuttd
Tf5wazlK7mi+573PStVNnD/moSL7M1YluEVp5D9l6MOFlzKu9TEonLijax55LIxmXC30a3wZ95Rc
6CECrNasFjAvrtiYcAwVd/RDSnbOUiMabQl9PrQj5ASQ2BKCaHGlTJcvStb+aFKFbZtaqq/ZZJtG
//rD3ja+9/VX37TwXtsd8N/eYLMftbDb8M6mTT5KnPzRazeREX7A5qqfs0Ex1PP5RTGGZxp0hX/9
ZAZYla1xR34VKXgGm8jJH/9Yuq9gY1ctV3VG+f4KnYR0RH+j3ujGPwYNuB5myoU4L5+wQ+QULCYN
tF/2fulUQVotMl2zhadm7cB1rX9OLak6EJuSgk+29y6oGXWQjvDDZciIw1igvyI86bE89+yxfacR
f9UXpOkwk4Vm9dn93mRCkyA7BluKiligt6HapVEs7EW65Ybj3mD4M804/RRC5VC5p9kvGpBEKdSW
UtCB26swekyVzVMcWVwOkEQ+MlhgLQFUzwnsZ18wVnD+8eO3csdt16OA0LIRDCq6p7LsUFngENQP
9d/xwPeoknk7kpWpxykFKrDMMOzKQ8ZecIfoAe9a/sVrhI4ZzGPrrFN85nkPLaDGInWwyEueWkgL
v8qt9YsDhzZEd892+kURWc35qf5OKrxHAl687rDDNsaNpQ9aDVHyphy6OSqI7NhgrmdejWD06HQD
/tcY3Dn/JsbjR5xpMe/aV/87K4Mp1T/qLU6A/FmzEyTFlht8R5Oyxx0UiEUJPKnIWUrOdeWu2mEd
VkT1uR0FrYNMrovkv6BRswmoZcY5d2bTZNXeJpM0xOWvQqWJpJFUi8wC4pqkYVwiIbM6ynHbq0H6
4ovaBacTbCK8+KlG40Wyl+PtBN9mcZrNzfi0kXCDPSnHMPvj5NnvhEvbZygtndWMhS8yiuevQw4z
hYlBNrWWudsaOXdZ8rl+dcsV3wT+8EBfPZGnP5Ny1uh451b1WVs08jgdV7ZJWKZdvrZtLcFfY37k
35mZPLnQ9e64ZMjN9X26Q4WiEvDz5pOE26M9otC0tbviNNMn31HAqDs/87tHr8H2qDRApriaKVeM
CX6DvQ9VN5/L20SQj3iqi4Kw4TsPXvc2MMfjUncmuVRASVifFbERbG1KyobyUInCCWnlSsXeIS2f
gLE5ZSuxU9/YTQU65AVl5Mk1QnCHGDNVkAhX7+EGyiNhY3oau2rByASYUHcjoe6nE63ocIGIdXy/
+bTwdkLtNHUReWOpgQu2DlkgmfmgMVrdrQDE62w/5pW7JLqRzckkFkmXnxl+azFhcEQuQOxl2DUD
ooperX1GNK/Ttey8sGEFDsNqaLbNrr+vydpTOFW3JM/TRrABY5CvQ+flNQbuQK3z3ULtP1LoA6It
tsOVfno5Miceed2qQuzRudL0RTco0zH3/fBDbDswG5Oscp0Nuc3vSTuBciyoLbYMtGNeV8AsRx9t
4/Lpx9ITlKSPRcA8NW++BwMjlB45bwxWAu0nGglXYZbBcGRMLzqHUblDGyMZDVT1YJwx5NSF12fM
q1nw8tP8gPOuQ1wrYoow3ep9heSwrZQu3OGAGxupTJY7xwPThvrFbdY23G8MFuAw4FgHlXOtp3J5
Ytw22bp+gtjybl2sUmNk4f2u9u0uQyann68kY1tU7NkQh01/clgE9B2rcLV+v6i/qGDJsClMOt0z
Hg81SbjKVH7cneodSRWSXAv120eNiZjEHQTZoJSePFmzDKEOCfngazuwaZ6rD4ZHUJCRPS4a58gt
sPY1YEP9J6YlIKgIWJFrqQQYpT0vrj42TedBK3Smqi2poWvs//8wgM+m6AyvANNkLVSCEgtBpE4V
Te3EZc/mYHz//k1xzb4wMS2/gKnFvYpo23NtvBkczPP8n4jbvMUtYdNdJThvQ21qaJRNfB/Q/NKO
cYGA/dn9RCN+WpddEYkVwiqL9ruGAjG562OUpqZMnS8kg4OSvHWk/zwq2OkaHlnnD/ApuahkU3xD
qSO0ngxmMoE7+wSoC/Ji6W+ovvFP+k7vzfN/GR1gzXnDvHJF7+UxHmY1JGN/AYPcUKX9fdMWcxsQ
mB05nLA9BWHEqbWPDhTMlL0a6DcacihZ7/ywaKmVpLNAKaYrzYzeiPWevCC4xdHZ5EKJJRLO/Xox
rqTlDNdUOOFtAuQAGahCvlP/tRlRf+4EqTQhrYdHRC3Abl6VOBYYy/6/pt8vZy+0DKdNv649buh7
CdSJQ93+t9rKEgsUbfqs7iPrSLhl2Ft76x3XeXSt5JNDag6gYNn1Bev1sJj1dcg565yFUJ4trHMI
bHxG7qNne47atcjFot3n9jdqvfixBxrPwyfj52fGJTHFNZMg6fvaBY8Jvn+3XqahJV1jmZMKsYfV
Sq42UbcpL7QUG/A7bJfz0OU5vRJiCsCVcMngZUwA5o4v5yZijdRCDSUHIEfNN4Yoi+C45q5xWzIu
hMAUXehHBta4YnaePMpMs3I2JQfLCfr30HBgik1Dp/PMxBig0Zzn3gt9beaVMVYXwbG1sCR0YwBE
3mDXhZgUzYthTbPWk0cfnOyrq4LIHXAKLe0aO5jPur+i6K2JmmXzesGctVNLBoA0jUH3E6Wr/jIB
A8yokJL8t1WZceJq7i4feJTrYqhtffDXT7DlnlWI0uxHZJlleFx9Ubw91YuUhxK+scwmUSVgc/ai
1LZdI+X01ENsegLPoUqMDqr1I6L2JwWW1kKost/4fDhTX1eXA7JwEZKeUHDSX3PWtpNbIVtaAhQ4
Fiwm3TFM2uchhAlaIeHiRVb0RRW43eNUUVCHmyr7YPqE09QreA5cYf/j+mRcIPyVe7Tal5rZR+F3
BnkcfSz1PkMa6Fo/NX2bigokXAiH4f+/1MEvtOhrBJRB7dcCCjMA8CzoIuY2hP8ZJJTxOleCw3az
2KH1sLaS9RQBz6hMofQWK/BxpDJZgKGQ/JcivUP2I6d/p/ecMFuPeIPBRo4oBVLySDGGpyF6Yn1N
SR8jTNDv74DIPS0Fdw25KXRyzjaoOKH+axm1KdnR0YVHW0ygQjbUD3xt52XZq76rLPHIzTe0lp9F
W/dkMpGGuQhF1N5zVkJ9xZftbDSLSCT6C7BgAVofd+VKvG+BVllxJsayeRI8p4brAEbHQ9AjdyOp
8reVMX+w/zcsjzWn4YtVk9eRveTIR4Wz6I66Zi5w89RWM2vHNq0XTT/puHj7H/7/7jBQ3kYX361X
r2Un65pWguIPBBY8xxu4yWQbcfDpJpKanue3tL3H4WgsvNvBzlxl2KpOmb2Xz+ugUTulfHAYqL2L
XgGuw2rhdyjzqaokcacDggFrMYIFjBhOEeMuSRb2lDZwrT5VGVP2SuhLa5l9QJ06MG1msNpR8f2h
SeAdBuZSoMo+sk0LYPiafRkQvU92V15rsc7xOMittc2KLkFB9mEVNW/Vu4r6M1BSp44V+omWBFqI
tE9d8d1Z3C1JYRQJb+TuQ6q4iTNgNMhctjB5mnby9L5romDAHPSmkYSBv5nhEqUGiH2yzOCIPnjC
mHpjcaLKnw46+W3xYfREhAB5wMFVnSDkhwNUFKISkZsMtnJR2MkZK7CJs/9KxkoVERD6ABAjldBA
/4kvuuXcHy1zELrzvJsPM1P3Gky4mU0HEUcGclSkWP+w2dAh6HTMhGg78HNpibu16HmU9258wq6K
NpWJOTBKgiYJAp6UEuWFaSlJpL35AATTin3aLtu4r1UXEYPEffzSilllFqqAq3Etc/CLT2p5stuy
PnwPuUOPaaEc8bZMbDbuF0xlitDGI5BdLKaKFjfyWxeuuPKPIJJn+yh9wgljzjSJ+kDam40+zifz
C86x5Tg4Rl2ZVOXyIO4c269t4x8UDMlIIUkSVsjH2Ofopwxch5mJBQDRf+ol9hAe9ITYv+lN2eGD
WuKHFXG6GT3hhZ9Fli0/CPWnBNZTJAHqk8ZL29JvoTVXj36QNqALnr7wPkEvqf1J+1RLe8ro+4Go
EMG2rjiI070+coI1QxWowJPUkbV8jn0C0DD6m1wmT92yMnqwUsaUatWE06IK/p+nEo7lRJqSV/50
4BV0XG0N4D5xpxyayLTovsSht3ScnVbtFpnK8VAX6K+Wi1gEJkj0pdysjBlBZaiXOErV/XthCJZ6
HbvE0qqUT6wWWRP3PLWx1Vh3AtZe4vv2ME1SHYwweyXpTnWFa4E5ayrjrO3xkrXCffV7dkIzoBxG
kTLPN1tpEVw9BKsuxJVQNFdEr7A8z8qANivIBD66/D7kn3E2JSBEeHlGOm37xN9ldz0yS6TcTyVP
1CvtNstDRr/Ot5c4g18VYNEceHABRPzg8mm6KxSFRImuWfNOeNq79E8b6bPdHxxP/9hBZWN6/RQW
55I9Cg4CN+Y563T/XXwUvypxA+u5kcGJCttL2x1cKKoBjcboiLrYOv5bGWBx7DOfrExDtDMrKfyp
MbopWODTqrpeT3tCh4y8/UE1CeC9PrLYRRtAcoUOuJ2AV+w1ERqj4t9hNFBrvwYtgnIcRwgQtczb
M8gZaJrVXWGj56P2nBj3jeQoEvutOqTsh2YfThQVam24GSKRhnlrH2Zjex7DKzXUj2YxN5SF7fzI
yq2NFjqJSUmQshGG2aqLKhCGjDJgSZ5tSYZxY/+WWDnKib8H5H678yOAIV9R9bBAAH7uVJc6pLw7
evGA+Er65+OUtOaXG84aUmK2iie2m7k6JgjwkBtjlGnXSUq8l0VuHHjyTZR6ZA8jFVV2uI7qvdmo
BUzxplHNe+9AlcFmJ7PgQ34HMZ6ufUkSJMWHFoKgWChfReKbUHAuHVH8qe6xCJ2zujLCs1FvT86i
zueEPR6rQCWbV76FE584UsB5wEGgQ/2qPx4TvRaNwVOWKGDFAk6ba+HSt45XtHexdQ6t1ICtRaI1
mQb6W+mJgVgU5EoR4JG/5o5xIfYN0HnpXJ8oCvQ53sCb+/Rit+of4e/3Ihffyeaxv/GfCTfmlOxX
gp+Y/PJinyyMJDJd/Aab5L9o0tHPzo7CpeagVievALx8M0ivCBqXmZw1Mxe2DwXqou+BTuqoP1nU
7ogj7UB+mNLV0coFfRseMZXnHp7zXiUFI2l094cmiiBsUnismnrU6eGsakngu40VCGZ++e76tA3S
9JrewMnxWqNq4A+Hu6ar96VxyK9cGexUug2fk3pJfDUy5nRPktmTvaZ9cVOE7NRyUJEsl/3xK3Cu
Tq2FNDqcLjZUu1CYQt+j6diMLMmPxvspAeLHCa/c0y+ndzZrBPYHpBRfnKliXxtSBf90z1r2LWxz
G2mGOi0Zra4ujSfUoE7aLVlKBakSLQfKsePOj+4sECqgLVwUkGdikj9fikcp6Xs1tX+bMKzDwOzZ
ZGjulMleA/17PCsmSeKtSjgtaNy/JMMj7FhkrEUa7JrLCZJKnGG8kwiAupdmpfD8mtdB8MfAQcT3
NoLS/OBBCnA83nAFfVDVSeieiyCiMiG14zEr3uwBE2eb29c/UmbY/gQGbTa64BF11gjmVVjOqcT6
+BT1HBSa4CHIvi3lRJzcVDjTHPK9khyrj0ZTYXlSsP6EZepnEJtGv8nA5oS9jyXxBSWkzu4IaXB8
hAzRBbGXlFAtfm+yPh66XKzVqh2b0sJ3HglovH6/nOrETYHc3WMTjHkr8Gp5hlKy+fnRlbqIv/jh
vfRumJYZsvZX2U/gMWiik0ooSSeWdYFPTcXkMi7EsiVQrKiwLfl5DiKM81LIZnYFE6wXNFKaveSZ
sqcFxAoEh+9ZLy7fZGhQ44WfzdvM38AtJlezc+vp6ocD0zhcpwiKqCrALFH4Y6h+20nXd3WByDtE
TCKj8jq1VtNIrhKx8emicdQTWGAu+Fmck6NYwSeMBfihRLPyQTSlb9f9Cdq/0afg5iqqhVbMfvP3
shGZodxIByLIhDIsx9N11zRXir6j19HhpkOJeTD3vxC65dK+H5+mCLFuv94oG8gwmvaomEtK2q1R
swc7pkR2RWybQ0OrvsuO/N349e4ZY4x1AHX/rsQ1svITTI+lGmgNQCYOUsaxG/vhNLnh8xpzoNe9
pfFg3aBmc5R2+N/iYdHnGICr4dG5om8h3Tjhbslmd7OblDZCuZfQsZyUoRpFwdNPr+HXtK1JaLUc
RiNi90jLeJ2agB2v4HPqjx+2+576VwKdyytrhXSRkMTz5FOJGPODa1qTsmALu74QrAJBLNIIrG+Y
9oYfQMGp8F5KYJLUK3K43+oxy3g382gUo7rlGWzsDtrCEHdRXEPV/EvxV7ssmkyiuVmgsPK5BN2q
j2ZHfHZk6AloPVAJWr6l4x3QBWVYWSuG/G2XgsQ/3o2369vovCW4ehgqiht8cnCMpDu26clNLd0h
i5nZrHhWgJn7DCKfc3HG+HnCcn+Jesj+jiU7QUKltAnhn8wf/4MeudJ4aTEdYkOI86zv/Cb5ZET/
qK3hB1P1HAlfZnNhp3fYMugt76N3fx4Yrh/nWMxKerSWvthsRiPFA76v85GwcqlILwleKKJGAI6N
o3dCP3ZJC+Fn0j9J/bjfVR8/iw8DY6Eq4NREFRU6iUTIR1EvaVMYOXij6aFICs8m6WrJiNesY1GV
Ai5RVJ8qPPKjqXvEXOR2+e+ybN69SJWbUUyOjv2POiP89J1cmPoj7K2eFBPsOpVHPkvJWtvKcqu1
dASkH1cx6y6xc0GiON2TgS+zSOXAxrcWscdZNp0bDv3nXj5SbCIAHypqhYjQihpG/mUErbcdr9Lf
YpbcsWCbfDM2/ZYQMPjUnFNIJj+gVhyaO50Zurv1RE7pho+rvNSKOhsPquiGFCUDJxwrwpOBFB3T
Va0pyt+fJcQjGUOD5QJsEfXNKk2iVIyOAYy+GRj+2n383UExtIVBAeDWZ8wphOIOWBRRb3IavCOq
MTCa8JQHwb0L/WxgMjQ/5ntQSVZaKb5C9Q085MrMR3uQ7+TKFVFzB7OMqI+2yuBd4O4k92qQfWSl
ZTUYZWfhD6YYnuSvuKezVfuX7f2/sduPy3gxgch31kniTaM+H6zD4jiALgZ5BPDQBVo4xj8PkPln
dQhrF0IMfPjrQmCNZWLP3SXuqmodIQ9KVVVo+RkxKM/jLmvXSy2XxgtN7+Zie1D5m0E6bEYiPwjz
NJ7aLZGnb++8W8nZpIAGhYap2+B6FOTBPk7swkFospTZN9LV7+q0R/IYDaUs1KaqaFLYFr+K6xY4
qMfgSJUAuFlXd5+LLqZJMTjIqBPs1x1g7CWWP5GRa1ne0vuptd4i4+PPrg4F23OGSfNgdTsOA5Zf
WU0QVCdY0OjlNq9rHkV42PRWaTXzzgiYkNfvyM4WhCqLvNPfi6TGFV34el5deGK46YdjIfJRzFap
SS0aU06KF8K8sOAigMRtUj+s2e8uH8x4nyKTjuqAYSaxOBji5yrFJE3Q0+ETXGGs25ShI6g/d83i
5uH494E1KIwQu39vxuWNjUk81m6GAs/k1wKo7qMRvjrpyAyufO4P/bXvHCxh5nIAF6M/GeJs+yDu
u0v+CWt8v+Y198AhOu4+G8uAhYtyq+smZNrrMmrr6Zfil5q+/OE62EmNSpfQPbdTY2xd3RU92JRx
+v1BYUFX8pkGOFTfkwrpukwKaByX+sjINThaAgaF5HivY50ORbtzavK+xwuD5Z51aNmH+UrINSJx
TwRokiQkasZy+0yHydrhhVsM+3qQeIshcmmkZPpgYd8cBKqdX3ifs39J8QM8g0G/Y20DANMJvGas
GdG7KTXQrrgKj+9TstsVXpFL/o9yUDZTV+fWBHpAF0uEuy4+rtPuyz5HDz0m4cItjMcqQLTiBH1N
EU9GYHr5IiFEedLfCsZAsbEZl6Pgr6IKJY1RktjCOgg1y60TIGgY8gNCLjMUFQ3ZlDoinEpfr2M0
3KLC59og6r0gbTwzTG6mAJuDXDj+UjBDS/X1rj34cC7PDzrjzUmu7zpXbpskQ8FSQuDM9FuHNj6x
RIEupmp6uQR64tQUD22NUKROUeTyzinKnfr6aWXHiePLnck1SLcsqLHybDRI1j9yywT/9yxjLXR6
+gbv4nj0cADs7EqWPuheIfTO6q0FMyMnMTUnzOSsjufLZxIA5y7Rew39CveV0nkEX0rWEe5jP5p6
iDCoSZTofHNDN0fLxd7xU2q8TNdWhNPdsioWdfatXC26qEtjt3wBsfUlGafWv3RcCIl4Ajja1dH/
xlZETCIjoi98oC+vkg/JCxZvmRePGl0dsKI1SGI5q/CE4R/kI3cJP+iRVNt8tB7IbgbXXK/4SGIx
ZbJ24z7kaiPfKvxY9WOfL20r4Jz6Pe5XCPeTu+AxTyZpQexapt8hQSlq/2XuCTIvCYIKBiLknpYZ
mUPFbkANrR1hSmSV4xE90SaQXv4Noei+v8FHTlk6tYQIIfh5OKQna2zdZbuBZBQi4W+hRQJvtzBQ
1Uho3QctqyGLSmPJWvu3YgPbViembI2y40NcVEu9hDAY/FRrunV5arrQVwNcP+DEIqlynwbt3+D8
ujwqVInLqr1mgT5OT2E5UI2tC5cJqlhK2cWgwL8YPIpCglYim94iCYWp8U07IPnLxdNBNNtPg+zp
SjsIbrxfLjYpW9X6HU+d/kXI/dB5E8PUdprSJxD9ewt6nX8YJ5zffReaS9KtSafgOENtJyRf4auq
kXdQbw7LyiNRgjrBfOv0JCKHSXrmwBEZCn+Yr2Q2D7KuM0DoXEew1x3jcVw5Cy4Pg9u6f8ISVCLY
mSdgaTpIEfpPC9P4KMF65xjl1t1+JgKgBRUt/m2UTTCcciI8MR92WVH+V64LlxmGB1QqrvmiGFAQ
11mP74F5tWgZo+GjtGogjgyRXTpqRXjC86T5FncHTLt+3JGLpASJCQ3UkSC07JwwLPwWBF/tsaCa
vBTGmsq/ZZ2PJonKpRR7EAGvGnz3Tw45dM7rT+TvC+6v9vp6b67Wd220DiyFa+gHck/Wh0Pr4JKl
Kcd/fYvMOVd5quZj3gEKHAGGKaL4/ccAp0Dt8j223Jg9JGj3zWCKHR7SVs2lD3ANNl9GSeNcZTcz
H0Y+CZ/Av8iRwcvKc45xQuJBz0Z0hiRroEpV+fX3cCYj8hla122rNf78RRreKGm/vDCbla3qQSap
QBjYaJBiWGXw41lP9KJ1s440Fr1JADz9R6+R+/ybdZOKD3QihC9UW4/jGOOebkcb/9gPi2EuChDV
Roj70tDfBgwOQ3NJ3/4xRslmhoz2GeYrIEf90h6BSWy61eKuiwPTBwCCI+LNoFLR7rtJS1xR+uJU
76zzmH+l9VgEGg9mZF6wwcOVOAI64KxqH1c+iJslAn0VKcDc+iK2ZXCRvF2ftkLvyGghcILZ54ne
8hoZPWzGmFrYcsOfjhPSMVqH7ib7mhQjdsAFssIqR+w1IAM0Z3/QlpfmUWPaqHr5dJz6Wqbi4sGf
BTZDEfXSXo5NNppP8B1p94hapzOOhf835/BXmxql4HW1qjMBlhDLqC7gdx4blxDrqP5YNNaoo7pP
tG3auJfcXHCHKuxVt79W1ts1yaqjMoO3YPAIEmFWns7khtnhZCiHGhqrvG95OJjrAKGZawmNG5nC
AUJ3VRAEvV7H7WS6aBTExrnf2IdUIvECDjGVwFNM5Jyz4HoXckEmV6g2CzY2T12fabjOpdql4rZM
yHAF9rcndYVTJRmOOkx4b/rhmptC4TQHa0Mu+XqdWGSVLoCEjx2PT7yW2Q0nIl+uePdUezt8hDZA
BYfl3GkNjunJ7MC/+CHpSZXbHkdZmPBivBwYgqNRXdFmp+GlxDZnKOsSTNnEdkQC11i/cgngERUG
uBilKPMjMNtzoMeyvB76X0LCzSfKi4WMEQaJ4q+thjtVtXttfyFMJm7mTchnke21pDupmkLe0OEH
9APZvKgV+acGJpopwjqVVGkfMkXl0njmJTl03NNwmtbc0nuGkAPAxIYnC9Lj3RL0bJDl+pe726Zn
CYyB4uvQdvliAyhmz2xwhmWrcxWdnoURjzHxnFslBjM3SfFwo/ldwke9O6v5+9Fj0EHqvbnNFsu0
B1JJn/MsTb1BAmERCbJ34ddacj2lN9aQZwd12zc5o7ZLTGeMlofKQrVebbFuf2AIcAWs9OTxqDGx
XrN5cQ5W52uhmVeTuqwjhnwb506wYGZE9FLMIGE40cJ6HizVNYGubxAe3A2K4gIjuunOomc2WOj+
lPp0OEAQo/WOfFNOsXmDcIJtv6JJdCewIdSpjqkFSqEKicdMKWEO3H3uizRIakDY6Jhl4vaVjyhu
/L6voNHe/j5EOzeTFQIpvVb3ePFWLwKJb0Vf7EqTdWYco9jNnf5HopGm4YJJnamv8kAiJ/jxQuns
Q1oqhRfaGqfnLz7LSdUyvqBTDxlAkgJLPybf9j7Uq8sQ8FbakTfB/j/nm7gdEImJ0n4xpODMAtq/
32KY8wXSvjIQ1wtkizywKZ3HZXuI+UN5puC0Nmoq2lQj+luwycds7BdeH8PNkQlD9oX+pvFAf9Ua
jS5sQcbIvryvPLAiKCdfc052a59MQoVxi01vut+Lh4ywERKTADnb2cnjA7um4t1I9KmydlDWa+TJ
RocZTeP1uI/Ts+WKKTqQ+T47fpbhcebuhfNKPqmqCU7QKQ0NVwLW3CusXZHxEqmY5Tk6AetDg9VS
AOg0NbPVbSNmvhpb8JfZUZqHEdRSkSTRfnjegq20YuSrKFNxS5oUvGA9yhjJCv5iwEn+P2rD7vWU
2Iy232gjmgbGiiye5TGU4XNbc4ZgJFzJhza59anLl49RZm5ffVc9Z1Z1ody2RMTJNY7j8HJC1wEU
tfViGh396fSTcjkz8y37b2yDZpJrpOmlbs03r4x8j/u0r/+XfeKIDAQ8P4ZugBzxJ3sqPUM3VeL9
aZ6jW1IqZXSR5T4aOK9W6ANxdB/41Wq7cFX5BYo6J/6e+uUaCCwTtuaHW3L+qZbEU+WSmZ9CuNbR
lSq+LX7i7DvEbo4l0EbD04Z2Rd1rQ2DMUrqck8AP/vqGSVRf2rk3Ed+x8jca3oRlrb3pW+xkchZL
/5HM34y88qjgYbU75eaklaqsIDr12fSHjIN88EoPMkkr20pmtho9+2X/pHy/cBJdCcUYy0mkxp6l
I5MlAXtZ/OmxZIdRoammva+WIIkMGk7OYXMU+UACsZDfS4pDGTiB+y/o5hD6gYbO7zE4aR2ZkbUF
JGbVnwIijOmPgB3UD/ftUlWXvZC5iECFp8gcgJ+EYZxY02CPxd/NIpZGT0U/GsZbNEuQpM2Z+bJC
ZttAV7tIOu8tIE5EvsbJlR9OXqgoNbaHpUGwA1CNBEXgCc0aP/AjoB7AZMgZWmmyMtlZB7SdWRcL
FHGQ6JxxhOXIJWttS3Wb/hyTw0C1SV1tYj5XzYGhuVeGWc06sOhyT17PpAiTYF/RUoYlCJ1MhxDP
Duato96ZdhWBTOvfz+DqAxY0XnMn9+0SfVq/LnaFJvEGqLaQIS63NLiFfX1IY9Oxw/aofb8qajSu
w9i6SzSoIRDRjW+RZQz/AFcDTF3p+s0o2gqSTWFCxHLP6mo1icXI7hviep/B17XAEc4hv2osRy9r
Wv2YaxdJddNvd1yaHm60AzDmvxOCOI06tmSillZffjowXD7ak2OJeab64Cjn5/Y95ltzL68lMDxR
2S3OuSCAmxUWUr7debYUiPVPNIcBycQmpt57HtzttClhjKKtLoN3srwGXCz/n4+hk4ufbfVVsUwc
Rz+lZVsG+jOPLL9v1eWhrOwDrSHh/v+rB0ZXXnE3isnYDvhUGXLbfmU8HVpNib/XOmF4B/3+voJD
O24r2lXFWTQdSRLOXR+32GRXCJAT6TjtzlBRXU9ldYeUYPIdYHg7o63OH1Edup813vsWSithOUBH
iib+TU9nxhwCZm8A0XmT8Qc6atkqSU/d0PbKnku0z/SxFl5YLuMj+CjbJoDGvuvnPzYMnm/Y86yp
0WT8nsLy4DkHYuRXtjALRksfLFt2SiunlY2H8bEttFJChDOND+iS2SMVo2sJqwZWCPNDG5EwwHfv
JYbAMLSidrbSh4SQL9diXX+SdywS1k6k8OmjqwS6lS9/NLqTGpFKrkMRLX/h1ozr2z29WDgDOQiE
qM/U/M69p7T4GtlvzAsEZciFmbFpDyALzXWLE7ETkq+NYth6eOuv/IFX8UxuQ7K3qGpO3rDzYHvM
9cAXsqV0oV+Y4RVfcHc3Q/Kbxhfo9aU8Z7I344+oq7XOGmXbtfi6Jnz2y/V9Y4ASWIrnT81HzSH/
yGwSiINoWKlAteQGGBUorDy5cD4Oexwe2A87uBbvW7WXD7D5eiQlC7oLtHoJDxU4ZV/EijJRWH/s
ed7pNosdgtPfGX8Qv/H7icZrahvs19g0I4vJND94my1+mFUR/3bbA3wRhGZIhOgI/9CM/opcGoWS
wqC09i84juS5HPxGSGE5Z1iTvbrwKr95vVlEWMQc4RLxf5JSpUjZMmgRACnXjfQdQZi7ThrKhqLV
klR4VC9+PzgFbv66RIta3y6iIukU1b9VVFCY54SZLqXcP2c4lYVCUHI7J0YiQ58jvkRn1mZvmAYV
xEc9bQc5Z3xOv3hVse3HZq2oU5sfGVGaacw09c+eya3G1RiTvA8O+4zV5QLm0kNjtnoCxdd+mZFe
FkYRKMlFq+WWajqn9knV1p5waNqrZFKaqVN4lMHPeaRG9Z+iBrC4yTUD4BZu7lE+/Yya3EoAyRp2
eh4O7sbGoycqvcNRUmR2fc2E5Sun9nviiDtZlOwkp8xk3I7JpSNfHXyWK/8jwm70kC2QyWd+8NUF
l4BW6U9nWB+kWMLaAvoUCWfbbZeb9gNJou3sPnwF8YiCsWsblQ0boYim3UGZ3iT0MCK7+4nQnVRP
TZ/El4znhEN+JbiT2xcZ6tQLiQZfqVdc+ZSwrqRtzv6PuI2M33F7PwxH789oXX/sesuspwvdsbHg
SAnKO7yaxCsjdrC9aT7LReSKkfhmtiWOyUyClzotd2FYP8bfOT8j6wZ8zVYnXegaLGuIbFadSnCR
/UAuqvpiXBjJH+laKXl4oNr/Gz1iEqM53QTF97olpWto4k0vSVAKKvbUz+uFHKUFiW6tZbAzvD+8
5B5j7wqljruRgzAyfmRwC9wMqKZTx5HxhDFCIGzDs8LYAL1FjdRdTbolxVTbmyRsYLSN/IeCsu/Y
YLwdqH0vyqVIF2SEngS3td4n4SNpK0WEwKbJYoVvo7DcSkElYP90jY4/Fuey+WEzGNXIeXd8ed9p
zZMXjpad2Avl13r5iY9bbVzOf3HYXmuYjIV8T3v9VzMSPDOdxRZNWEuZXOZXE0qN4CeOe7wgR9kN
bDG28rBz2rvPlXEuix4MgpgPo4rH09OOKHtnhVgyFusbmUVay2zy9Ay9cWlOvzN3LSQ1q+dcSbrU
zBjB3JXWm4q25QzaMsXN3Pnmn0IR5kxDepRbuGU+MgHoZ8sDR3ofLSEYDnr2JiGnmuN9bjWflXmf
fA5vmgXuLzC9PGgbdhXK0Vbj+0Qy0LBeh1D2Yp5Imq+Mu7A/2dfGSam0UD3Ijv31oe8uHYLFDnZH
Sv61x7BNKD1eaZ/1vkDLjrT8EyWutgMgmKTBtactmRPPsDRga/lvTzL01nhKjiwt68yVTeE/XLMZ
lXMSL+ypNlTr/dxLw494whq68jDgoapPvi2d61vbwEJ3ZO1NQ4h4C2DBUSfdwAYqG7PZ+uEjmTNL
aslnow9qGYv+wtnQt0AApAzGkjH/F7DrS0i5ztidl+Gr19nObCF0ibNGKj2cgHzXdHOmz/f3puoD
OdhaJAaAg8oH20SVsY1KlwX6QSk0xNXrr42hbt+GH2HIZpKsc5mF9Zcd/+ty/gMYUfcqd6D0O8xV
Tgf3GSdD/Z/ZqnBDjaF9TuPx56vpOVAIFN/XfmHckdP9JCPe55xP5TMlhPw6mXilM+WQEwn73u2x
Hp//ipQaOUohVDMrLROZGWw8xk/t2vIDObTudzBSgefLCciOEiG4DuAMuv9MMm1A41gaW6UdzBpv
QaYWFCO3fAQPyMkyh7Z/IlYAp/WXr8BpBizQA5dai+b0uudAYx1x78M0Zfb/98cbTcFmMNazwBfM
9rZYjKVg8zZzuzHKaGR0YQx9YbIdwM24+SctAAIn2OWM0PjambWQMTVr0pq1r63/vXP144ue9WAK
svPi38UQqPUJ7+cNg4/TXS+eWkZcdoWJsyS5pdN4fUgwYibu77L9BSAoAX/Esu6ViO9olse8lHsE
/0VqttWegYPAUh0Qjx4etZc8JYjQ7r9Z8/6iXyVtUMJ8FVrD0TvpfNjSd/y7hzDWAARjWC6Lc+MU
kFJvXCIPWSkF0Ij+YSovQSnVUdPmCIrx660iGAkr2pB+Tk3GPbPGJbYYc4CTvSpv40Ne86hiAKWK
KepCNJYs71OLH2hBQoZT1//OTqsVDjS/q0CKTM+iyfQIGhQhsXvuXsez+L9nGNqi1Q7jyY5mODnk
9ztG4t65cVzKzWW8Zb0tqNrQgQu4pjrV5fLJZeqzWKUp3e+Hfdkj1yzZl7ieAyT/N7hgZqrQTglN
PNmrVJ8NPe1nbiJYmFMAldaED+LkAy+bJOgAWJQQLL6XnIO8kQDu5kAFh29HkU+PYSTQylFkEWRq
ezhf7UC+LZ4o0HtSjOfFaQFNKtloswBH1h7kZfo3G01FB5Shsgk6cxgL0cjHJiPn3Xr1UpmfJvFG
QztXkQ3eXghwzhbgXBio6jPwNCsF/HlYLnFhD0ACMSaKNSg8GC0NCnHVTqyIqsqBHEOFSid+957s
aLI+DqZ4u0Ba3eRjDQCq6cInbJiwJImPuWCUxMAX5K/EvMjNLxjdHxIcqT9R2LPiCUVKzbehJAcY
fYye4mCJFLqzU2nc2GnGN/kl2bcxjPf20heHmubw+4jNLjSfH0Bb1Gek6qB/QkCIb2zibC703dzL
623Z1qZDoaaMQQ25Vi5hLEC1A9/gAIVOX6sMoXBsw3l9VaGvod5YOznMVucCxrFIryMAwNek6Suo
6fnkOOxzPjxEewH8koNUHyxY1M8PXAxbkpyQ3Qv0ldokLUBlvyKwYNVOWpcObNyJWKw3nNdfETX+
j8T+yt7L2bHtRkwDA4qmwXceee1X8jSlX3Ldt9Yo7SjVCgyMiXyjtKboY1vGNqGFn/xbmcI67HAa
R2MQXlk5lxEB8O/QGcQV6pxdJrKaS3oT4sTdDSupk3bldazrfQNDOGJM/nnRPU0R+czcetYqEPrB
UkOGOGxfe0NEr3QENUEwO4yinm8HkQc4SVQsZf571KsPkQy0MS71Ved/C6UcMysbd9/BAFZG6taj
iI1pOjn/dL1IUSjhccpa4c6LoT3PVVjOp7u20tTK7Ouhi80xn0dCg21q1WS4DYQvsMX906XeUN4n
L3VhSENKjBr5QoL0I96zh+p/lVg9mmb/uChSXoiwXcC7bJI5r9diTZGeCf1VJthe2Tggj6F8xTlb
j/RldHAEt21TBCbAdiml7rR2baonIfh3NlNUUatp4fs8js3S+dMacheV0Qiw1HnywYowswo3Rmw/
tR1wXwV831SH6SMziQG8f9pY4Svv0BEFEZw4zXCWuYThQT7wNDbXGxkLKzf3EYjesnJurBGqgCQQ
jKqDai9jOMtAEZhV18zfMyAW77SSt3uxqXhX7hnA9EnH5DMCsMDe/MSeft4EAz7hITVdB6981zep
WIK0WZjo/b7Wgug/88UL7tEE8GZPs3ImGD4Ikfkanq2g55JTAqQMAuqe1m3XDTZdbNFpkqLysmmh
i9Bpd8/WevxX64tYv3CG1uD2hsIkuIDkV7pPypmMbkxd3Lhk+laqunWSxbCdopfXr4Qb1ERsCalo
d3EJ6CIY2rS4r44ovEm0fJQW9vpWU4vgnXB3wkgnS04h+jPcENPDDMQOquTZ8l7ojGO/mUJwoqY4
XtYmXM4DNuZTDuJB9KUNNc7u27Q4STxmNicmhCThCtJ6aBuDuqAcPtMg9M9YlgirCRC2WgUkCFsT
PJNq66VFB4isUB5Ue4sNwHLYpisexLmIytKkGBmw71IV4S7mwy+E75IQuitDiwR/8N8Od0poMQX9
7anGTJVKBzeAsXVz6P7aqkGiGACNrds5LmTCrjM5lmHuKSKN1NlcE8xZXhPHpbozNdPqkXPQxeiY
P5jPBljj80LXrEGOC/kpYNIYkjpIsDFGkw8usxR+BZuVx0stBjClqSag2G5xYu7EBOCSmXhiRy5O
NzQiITInqsbrpUgOuFmxljbARe5loGshmxbFPJp74QaizSCaNlkClZ5ifQ+YmkHiKBmSSNb0MzDK
VzQTmGwa3aMvyb6TX3W0kzWIA7/Qqy3A7rE6l6wTj9w2dYQJiM6iqwS1EvrwT9fFX58qAF30Tx5W
C+M1wGwhLZcrgTMMCaxuIuvsbU4sd3bp5EnGuQJIGDsThVsIFDBAPkk08HhNUIgjqoQU8b22ND2A
Iqfkdjjv2KcdXlb3LpdKB+Qvuirot2wsOHMgm/XEckIKhyqj6/9XaLFH/XujViN/qqMqiLWktOwD
/Pz05CyEz4i0HShSFBC399WCbqSWWpq3Oc8qQ+Ygygo7eEw02tdFn7FeeVR5WfuEx9LcEtJHjP0W
Na/2V5f3oZBWd6Af8jFA33voLgAEPDM6KUj7vSwwohPp0XF6d9Nm6B/kigeq1+tQbURcxmrkqkVs
GrJPEUdpDyUB6TNrigjhI7m9P2GCOAdWuRga4GG44HylymQvXfMyZYyC65gZ0xF2J8Aqlvq6jssQ
HDORnixzfYHG7Iu4j6KhnADWuCjqYga9oe+ztrmuS48neq5qUg+WAiLaQ289Einjs1k/DFlUW1ZF
X4eg7VP68zlRpTnV28+ZRy6awuga/it/zf+B95hZthZQSPZkL8zUZe9A0liTsQxoVekpiw+kF/9W
qKCnqzBXGgOJ45q3jMWuoUV6W5VZFP+G/0lFUzXga8E1rLOR1W+h2fuPiriEEHtkEG+qCNEhMtJg
luyQ4jpy2CwI+4fT7GYUoVqvHUvWmkqH3+GbsvvL11nE9FeRCwIvYJY0vdHojMKD34pBoqHkBikT
WIS6OKXKwvlkdPDMHh39fst/px+KfS1oed0YX8LN9BsfYMwieD4IvpI808B2JC3OZnaytD3iccCr
IkvWDqZle2WzjVLB5pU9B3BfRVNe48lcdmqK/uzz3qZhLotKlVJi+ccB78Ck22BjsES+qQnNYfah
iyvxj0XgfUyhkSvZWstheMExpRIHkNbWG0NgTMf6C2QH+sGlV9tQgjLz53DlpESaP+YhQMgEcuA9
X9N6jek3Q0ISF3cdHL7hXiGR1GDHZT4u1diwaZ97Tn4uy80HA+uWyD3sFygbuaZLHmcUXtqhPE87
o6Prwwy79ING6m1uHaNYC1JT6TqrbQp5fux1MF8cngrQf0pQ8gscVjhDOMFg301X/qq6mtq7dRAL
+GvgaEoVJosLzN53FzR2ppviN7StJ68/UWLhmg07NAEk5/h0AADzjftCm4pnGQH3DKRlOSVvovmu
3wBgsNJLycaBGjX8W01kfTSAPYngYB9jtZBteMrWtRwt04RKsBkmSbokNmGLL8fMHAVXnDeuOvDW
lr1Kr0WcMfWWPs9bLyWBzjIR6ln8ueBVumvGDPGpuQASkOqxjp+e1sNOmaEgspjKjTmiwTsHinAA
OwZX3+Z7EXRzQucqwDXoiiaOCEBLBcvZuayS/J/ov/w7RGOoC1lkwJ9D/bw/69e6vRcRB3hi6HrN
aDMK64dtVdQAUIFqBYP/eht2YXRkWh4AeEurE71DYlVpCg/2uHvYXVSABjqepGWxFufcDT73DkIN
Ea7/6HORPdC6UrkOzyrZz7cazSoCVLyCZudGTjW34GnYJ8Wn5rO0Okwb3kfEt8SooDBgJpguCBc+
Z4IZBhe/w3K4PeFgTXus0XokMQS7N5FxDTZZFxPk7TaCdz/G/NGO4q2DZKxj+RX8JzI678wl3Nz9
p8212vxp3zeQcTh4XjNuoLoois5/Xp/46PvqlnTRTkEkHk0BmT9dyEsvmx8oNx1pvI9CDz1d9qiq
MYa0aDDG4OsnplehCVjcifzUPfOHqO+WbM/38RoqEe2dh3soAfL6XGBgFdFfnksWejvSMVICJo2h
vYasXc4DKRuwkIZxnCXx13W02rV5iLu6MBGZwjKveQqPDdeNMAGsEjtZ0wFaf9V0g6pPqx7fngZ/
7RRjdBOLnNFQQozdzihRWqYo0qJcszwRWprZ+RYEivg5xs8ZLRJZADsznsSEZZmINf9yqmLDjDV0
uxzWQ/kVeMfJI7wb6CZtdBPA9TTm4GCIzmFfCUIpslwRKnKq5jowvOV/OAA/d3ycRLfWs60uOfft
qD43Y3NANIMLwjKHgMTniMIdinZmE6/ijr+KQ9UDlhB7xTL+AvsifOVCt64daECazSFxt7a589SK
Uc1uQNjoEei4rhN4xeLmxUzqzY31I7J6a8wnUaeCInEnoxlN5/WzkgWQOfEvXC5Tf1Irbpu8U3v1
SfA1suh1iKf0E/kYM0/VER0YkK7qRsLWjpiJfkvhOPpoONGlPf56LljVV/emM905cB1rkQrRWpm8
UuzWPUo6Tk3VTNtH/7jU5x3HjASJqh2A2NmsRTXcLswtHqkNgA9BTfNfIXMo4CmR0rCo4Z57e4kh
1bbT57KAY+FMSRvy7qz6JwLdMFgcB2AoLAWLINe3zxwlaXQuSpvWnnio47TFe8OOZY0l40H9YTE6
XGeyAXlVFF3Pyj4T8U4od1nRAmndfni4De4msa4cc38ZZLphcN6hzK7g4DvA0mAIbQNKgS6eUlNw
BXSlUyFlznaiSvXltDWnO7BvpXijPnKZoA53KBPyv2yKO/bYseslSWGYHv0bUZgEWiFMME3OEi5k
T7zDBF8IQadgiO/ntb9B8TnZayZofwxUGX430JnsHE3e1EmDyN1la46+L0jyViDxqjR33JlszP6H
vWCzyGip6+BgHRZ+y+sNu0GRFkLHSm2B0fDxgTkTB/DL9E4NrbNwXqSGvKc5Jz81xQDbRdw4QRNT
Zo42yLEf4Sgyy/iRmxjw5H11CYn8hQvUUaNeA8vMgm1XLFlsVBrrR1qWDfw0a0Vjdo/pVrCpd62r
P5qfPVdYWBa2bNwqEww+19401lhQm1PCBlQz27Ybw+bQGuv2daEcUAQGxLMxRqQ3XvtxxFQAy7K8
vbOQPtgb2+Bw2Lzo2lt75MqWoSYRfaBUbo95NlmXsEo9oSYeJaEpdH+WtXxHkP++96ISXeM2PqOU
jtEnfbXglW0vbI7itMPMKm4naNNWzlGac6eYU6c5H1FcKacZVkOVooTr0dvGWHEpZ08tQK3Cjxh9
ePpVxviM7mBd1twyiEUhk21SMENyvDF1MwiIVtZVtbo90TW9Sm6SnVhHuK0WIXCoyHxd20U+twAz
nQncI6UmjVbnSgNECxHIz5g/19PIvfs8JD3AzR4io5YkSqhZ71ucVcwcplsjCfcgieYl9Xr1caU9
CdsX4cU3Zi/ZonUB/kHjtVIlHWyynNKnQGdNKFrdQQfZKbfFJUVGM+OOUUqS1oeiUmqiIMybeS0u
BZdsfsvkgt9fuP7bSRJ5tO58fvTwA7P0sX6ZGapXdebm/Uda9mbKnlIn6Inwnz/3vfFNBLyS7Ytb
0OCdd7e+O34kgqHk/BrbPMPvruxEuphRjx44rQXz3JQerYyr604lDPfTh+7I6Nj7ZuvYS/dXYc8a
b3UKCEJ6/gDox7ibXlfiXMd9AqNSIehU/0bHrjMQNxIoBgw+gM7jZT2yzPj2+tul4MsnFgh3L5ZQ
bv1vMsbELQSniMKmwV9eq5q+HdLamaNuKbpclBHBHMeIVifNaAr+rEXCVckbbGYk3CE12ou1RPla
pHRE5emfpZq0SA+xQDDTeeyDzVKl5y8B09YXo8kY0wI8Gt1nuVNI0LVIwxfg/vz6g895btpl90vA
u8+rjDNlMfgHyxFssmYawQiDPRFAsMozhViAk3IfSrtxLaQfENFELxI+SXXXRyKtSy5684NgUCJ+
XEcJEYXgkvM3GjLuKFvY7R4Cwjb0fQCyQqUi1tXBdRHKg69kP0n0VBrfIcBbap9Om5rzH1xsURNG
N13YUxuiwpOxkTKQ042wQasYdRfjNRzePGHWFrBAxFzv4ZcmEsIIeiOWqWPFrnb98LPPPzs6wUrU
qwOMeB9C45DgtUzYLzZVbCh6mH+xLJqIqIMPLpK58Cej8WL0+R5wEyhNa2FpH5bK8dXOiNQBnhLE
Zt4+9rigMekS2eAO7gbHnDkcgOazF1uZ1VXTRoOJ68K04Y7oXu7H10Sfo5UP54K3V1j/ocfVFwnw
C/2mx2pnbMXo+K8Oq9HPr/xFTeIUgzo3CoPGuEUJsJs9xNJMWuF1vLfHQF2q9Ix6po5o36KUOuDP
WIYXmra0jyv3E0mPXlXWJqoApOX/ktJIL578UuAvhAZy39WTuSCgzWNV9GVBy/13BeGLvwpAlBIK
8JnLzUF3sXJhg1SoayguDTPj3LRiIHw2H7SeRxsPpnkZOx3ZFC5cGdLkK6Q8hTJfwr/G7WNaxdyF
SkdseBVKOhyJgP2GRNoeSJrHwVlRIF7lX/V3AA8gtNKQdQM9J9kv8hREZWqKDof3+aUgW/bcRMTT
yn8H0Pnyj17ZgiRLa5YEs4fTGy5ftmOJlA9H2tZecVtqTWH1stVSrj+aVBLkO2582B3F9VWiMMss
GWXw9rWSE//+vPwTbt/IU1JDr2CGwJG1Ou4e2ga/1pFE7Cz0i9GaNCV9QpQQv/w0nnvEnMHZo/ni
Gwr6W4xv301J9LBOWiJo72acN6AGhYFzDtiyw2a+1GNdi9sTojg5lLZjQvb0k9VXIjTgAgQPjy1i
TZINm7ZDxc5QQQCp1eDEtGp+blDeUNAEOkW1q3x5R6keXby+4kS0zLVZCqbyi0S2IZJOITVOiv8m
MiA6xXp66XTDlCR5kJpQwmMwW9LG5hk2eTvvFK8zHBMv86U1GqjB6M64EJ9UJmAmoXaiXYJQwsCR
rq+4PJim/gPl2HdRxqHn76q6JdB/IT4OOqdWwDqsuKbh+9udfRzWT05SSAfiJoLp4sMqa76jKNys
cvJ+keonltiIkMkA8VLkIzQfeGwNCBH5fBUzW2ONFw9AGD3l06MUeVt8nGEn1y48PgEVrBXGaBGb
9klBG1roTKjLxL918QZ8Fm5Sb1PkTLxgp2S70tOtRCDdcO/67FI+HDF7eBruLz60hmrkuPEqAyu0
vgBoW/bzrw5EtdmpKAVbNvIGlw0u99wtF30gDjAMUXcYHtTWjYNtD55shX3ev95bxG/XmKHMBiTT
2pBHFh4hsOgRkzkaLUpcmmSO4FGroN/zsYENjTVGGFTA9XuaRbP5ftQMcsrhKfJZWzEN8o8FgG6J
AplnypeWnKwTuW/eWNCNyQVRyuNnqvvH7oVmto11AGi7xsCFc2nWROOLca0cjAeVYMomL8/smqeB
cOeEi8qLwJzccpM4DZtqC8wdWpCBECXVX/qVqlrID3uxsSo/P0alfhD2PaHq7IfpibmjghtGcpue
PbWyBU5FUFmJnKFaagNo/1XRis7bacSuV0rMDRzrivumu+w24L/ZsHPyFabK8XEYEsmZVd5E39m3
pdjlkJPFK98tHeQn7JuK3reie5xlfKBsoMrL22dKxLQQsPYcxbNEYdWDncpRBb5Avu/1JyL/f0d8
l3n+I5el5y3Px/TvQalU2xJfdsEH+a5jtmY3jkmqI/pRayVHpsMUSvVsH7pqPSZ6o7sG3P8pC8UV
p+XN+PSDf+/jW4EVuC+dkv9k0SYPw8oGzcl2zNoM1HD1rgYIHSOQdCNFFiI+DCbyOicTdzlu9gDV
vjYROI4h27bvxrLpacpZB4L9eMqsr/MBD/+bDH5Smu5ktbvh16FBHFnwdkvOwPduZecLzSCn37H8
coO7MZdJ4rKrrxl4kkCg5QzPwV/TzAon7fKVp9yjNxvbxyEJUG96tj0695sIbRFxdsNtWcq2U77h
IAyL1/+ABW5vRtatn63M6dAS91lLQAlZlI0jSbehk5Fz/VIJ27Yf9HB/SvW4yfHlI6kVd9XevMtP
NY/GxnE+x4ynKRWZkmhKa+1MCIEkIfXVjDFmGPrJxJiaiFv37YZOrXKxQganHs3rEyueDxkFSHDW
tz9WtVZULG68ZZq6IXL2CZv3CAZC69RJ38iYIfQUIqOdpkdT9gXS8zAbtTSOm+dc6vK0Uk6zVoTU
+yvISLs0QTeiYRUH6JcShW99PnmxHx37tLpgaHwjWGTpLvLc/9HlAfqtDKwPVW5eMEtsNl5jbS9R
uF8JPSMvv+GSL5LgeqP1bI+y82Krr82OWDl3KQj78zUggekhldXepdCWFZLlrzDxK6vCRjrFj1td
tZUbbjZhbHKyJubV9jg13t0KWc1LqLg8NFZwTPaPXguB8e2KeiDpzlbWmCCcaHpSpQuwuu05X+v2
88CSWE+iXvbcG5NfjBlzHC8LUI0oigvhDK3ibUB6Azbd9JbvMz3mCya3vxqSx3/6zYOY+jmaSlYT
H905javu/Iw3en+10DTr1ES5fIb1esP06uTDbgN+6Qy/NAE+zIrOIHpA4BZKHSDU0mBlun2JSawZ
Kk8GpbWKLRcLHVc40UwffPHcRUS7skTsC59L+KIFTTZT6TNvzb/X9Ub4ae1Crn9TvZ4dGfC1qpQ7
VFzmqj+OHQSdbmQ8cclLcg9IcqcmQir94Xf8vXe6VyOyZJ47KCxzt4tIvnPvJ5ISyRVcgDaFNjeL
2qRVGRkmQKitd/A63DH9SDyO5UU/yb1N0Hlf28qLWYz6zAZSB6KsqJiJwrN5iS4If06SOlI1T+hl
kgCv9G4Q7psii6WXHOGdhWNEgOQqdA0lVld3A8dG03781uLsVSNwQm/p6UtO0NyZi2vl2I2qBjlU
ulc2d2r3kTGNzlH+AfxjwEXPXGHeL1BGe4Yx0JNqPsjAjwN6FAKQvqNe7Vgu9bzhLKMwDngC09hA
xhbkRHs9dh2kGAklb2XMXtU/GzAE9E9Z0Uu2cG3MZvherqEtMDIaUE9yXgEpiLNboZcWUBdqZ8Sy
dOwF43lY1fnId0SIOLwFPAxWypxC3SlveKzce3cUrNa3JmGz1zU/qb4fGWFX57KOUytBrWZykgsc
Q1zj8iw+fHnwqA3oehBgcyVZQ+1ZMhCMBAioQRA6wjJwXjPknV3AWiJS6xU3bs+3feKEAxC86CcD
WCmpVFeFDy3ak1S9TNLOASrAWqI0HpFSAqEOEjVLVviCPAtnR/JWCAtm+mWH3h6RoAZNqbZb4Czm
YryW39UnpOu6v7Ep/E8fCPg7gNZjVWbGIEw1nCzk7SxGByhHrY+uM/G5RCxRBAfmMAxYUpp1u6J3
R899JmXo9q3Jhg6G8OaMjs2UyZeW9jGg1NnKMcv2DMvMTGi7X+/iXQYgGQf++plxmdwKjT8mveqT
3vIGDltjqqtGtLBBLw9bzxNDGfYi2Ess31HRgeqlmzUsuyjzGMmeVdIH2ILlXvtyATWGq0R8eHNc
jCZ3pe7oCFyQ0iUr4haT/jl7VKUcfaLnxDWy+LB1v20J/VkokupgLn1T1uEWjR4cKliXIw68cZnR
uqAmdfQVdBOsxb5c3ltSZcP8qXdeqEAsx2j0DiRZJ90jZkAWS3apw+C6x/PY222uIAbWuOuvvhau
9iqzAZXOQGlNGH25kUORprEEQuaDlN3QcvOc+LWJtpyYp3zNzEY6fcx5jdQ1NPHBStadb4vzPmKX
8vZ911VjHI+9FGm0+ZDcFSzXmonmix7ou+ugKnvH8UexiGCBhbDgosonRvtuSBW2912OL3HUE80P
24Fg3R8avdgJInFtWTx/zg5VhmQr+0OBm30jDGRxo59HTN5jS5/O0Sex3vVJMdWTcKe4YAguRgeN
H6J7WjdjEgocnPFw+wQ0+kIXX7NQqimKLcAa3yMpfBrbE/2W9UEsKkeVLI3NY7GDPMBfZGDU0qZc
AGDfcnk4z+Kt4jbGS/oOL8PWMDJKoUgT5S17ty37xXA4wRxLAN3ICByzfNUQ4Ph93EfLHcOvoNy7
Uu49ByJIQfn33524gZCfUaOY2WHCS0Iz7HNq9hwoXZbifPcWhorNL0sI3r5FNny5XJMumLb5uWmS
zwB6esEJ91PHdTkDuhuYshUtqNRJAzIg5zpJ0TcqrcHLgAg8n75Ptl9CHx2jBpKX8Tq1pBI7Py+P
SbzL45q/HYOAtcKl+eXVZV/mN07MGbL7OpA9vQSaIos7Xvbm8/fMpYiNMoSmHjkqRTcqtlj7E1rD
s7lS+/ms4FAF3wyzZLxio7G1sntMaWLIRlKjFVhd0bktIlBy42tWK2IVm49EnqnYxvO+fOzIlhcQ
fj9mjMOkAge86kJob32pxyosfsTS7p0VqDIxeLEHwrAinezp6PnKlzSM5Rzan6EMRwWXF3wdARRe
LGQaKv3ZGsdo0Y2r9FJ3rMmqLMs1abMMn9p91pWxAEj3xDlYRpBvRdZYLrico0T0XGH7084pdXBR
nohmnrXojFLkWuQ0xKAO07OOqi1hi0UlZ6Voaa44ySkbeMAXP7RvJgPeUTJUijYzJeWZaxfy17gu
0/iFu4jkdvYfKi70qeXecM0sNZjuJ82AGdBWO8CtP9G3mtSMeT6YFpYdwgjb+GcarazQfZH1i4pf
ghtuSFEKGRFuSu+KNVVq+GmIAahTgwcAi4oBv6qhaP7ya9iNfjn3KqThSRCusBMoFI5KdxlTdIxS
UMr0kFfcOgGNQc28nLUSgxjuKkdxovaRh32yDMuuuJEQYucWHsN6IBnyFtX3atsNgotRSyssxJXn
vRQKv55x/shx/8vdEj2qZd+UTll45jlb5TcKW9tm7mAz/IEqbcz19zDa4uu7QBgJECF8y7epnbCc
DQDL5127vxZQczqFTH5FcQcQ6tSdL2ycjjOqSG6BpI8YH4VK6qkiaiQvdzKoLyLcuT+5bymzLsWY
8ZzHYBdF2+QayGJJw4srjbaleGSiG2tBmYP2P5A9YVxcJM0jpVuIxUdG54LeSEWXCtbhy98TC0wm
MQzgCfuy4rM95Llo1LwYRNBzXJrTmeeFp83fa8j9CNlXLxwKTACY6ZuPl/GS04zZ78RUYywMxSxK
gzxS7x3vl+ZkdCjZX7We9s2ydXz8MEgnGEDVYvuehYavUKkDkBlKQRNR+14zPTI5pRsDhhhMDkNU
zeJQ+3yFmopKLmSl/hJu/k/7J2mM8f9M4LCrRJGJUtM6m9ZkhIttn6ZEVzG4vbzvoScrQv2PK90F
Awd7JwHY+8vBOZs+ps5hd2W8HhUQZfzZdkmt39v8xCgV7YeG3iqySy2eJqTuJUnoJvmIHJEn9O4L
2gD9B1luJlsujraUDeT3YtP7JigRbymAI5RUCnVYP+NwtzshhInCi1KdS8RMC/LD2AM7qI0lQSsC
gEOB2kgkjydGGE0S30xba/JWOfHAIOBUcvmqCGkckdgQ1I7YaPWUcUa0gTpBxzqLPr1zeUyme0iD
LYv6d2ZdICrUxfaM5ILr/XBASIie4UtpF96dCH65K7S+s8zaz5b9r6IkT1wxzPb/hOaIGQWAH8NG
s34HZMg2CpqBXFDi7STLajILPnwpxtcDd45XnFrFd5yv/Pp769yAo8B9w5FCSfooWSvwTGBboq/w
h1HKQ49yoWkhzcEBKSBwvzVh6XFTHhoF5ojk1BbqbVtDInW8DTpPe13aVj1zVfxT8vhRTXkJObZe
+FmRMwZ4yN8arkvCdGlw8BjSTMDRl7lJKOaWnDG1jPqf28gHXii6WdlhTcIxT+SR+W+OA610SNrT
Gi7cWmC04168eRiET/No/C24p21S5Kq1TPZ2wH7pzqPbgn/Uev9uLoKM0hWhvA3wT+pnM8qNWWEN
hNGDjsz7/Lnvzdj37fxQu2Ig38ryZ1wIv43T+3t0wIMO7FnxQTsqwbUaPJrK/20a7ETeWcqX6I3k
gK8xn1746Hz6ySbyYXdTJvm2P9lNjouvaQ3LE950SKiWH/GVa+ZcI87pZGtnHK8LXeVquVNxFTsx
t5w0ikjuxtA0EqZYiedbbYZaPcnW4js9Hn1xVksB15q4xXomUn80j6UV2YgGqqpRnfwfqhoYTJo7
1jY24peZ28lV/Tf1e/RsC5vp/g9F5uyulE9zGkop/BDAFpqr+GBVI8dK4JQzvZCy1XVZ3D3ZcAaI
ucVBAu4sp/YAPIw3ZK1BSRqZKq3kzNLV2vQiwshRFt/ReG+UAZJhzE5Iopyj2ur9UqlJvoYVPvBW
eNh2fZX7x/BE/HPUdPq5DqodNGRx9WaFyFBT+J/7JdSB/8sGc72XfaUqTNEELTNmAbwFWfHXIsmh
rq8LCfYIASwZpqB9a4C8G8QbOFlgoTJfJWz3tMcy2CTaYxHObjeenPAcey1BA9jJTUDySIQc2ZCX
cC17+SD9381j+uligGEn9UwPQTNL7IrypUeCjcihkTOUcY1vh76huxvYIK8pnjJdy+FVjT5OEb1C
FMi7DoePBGT/NBCS2WBIe/PR3MKgs2Z7ntuXQZXdJaQvX61/Jk2UOVZCAcHzB2Yd/Dgv9U5igxCQ
HfU1OnmtlP0TNxrOUw+l/f2XJaUFujjUhhx0AhyAGNRLKaOMSopZrM6iDQSEkjxKT6hREPN4DbJo
f2gJfIfI3B9eT0OdbXSQ47BIHWcsLAg51qUcQ1E5ib5CaapU2GUg0JSCQL5xGRB4ZIaUDJwWPuU6
NRQtFr56ME7f2WkyJpqQDnHthR/ta23600AFutO/YtPLvi6XJ7NZ0fUg5uEDdajeyp5rwtzXnfPg
nH4kGzSTHX22NwmVWkvz0CnJgkfSYlXfV70LOH8SrAzGQ9cN/q+cVu0h5r67kijDM7JiRYncGiBG
971dShvM3wIav2hohUS3sVOR9dLQ3Atr2619op1MdRuQWaYh3HRMtBMEvpCPXKPtAeH4cFpbvQk0
2xciVC99Wv01kCQdbdo2nWibkyEwNVXXQWYw3BfdXdVm6kJAwRDS9NgkJUurh0rfNxb40DY/WdqM
qw+YdzwtdM05j2y1QKYGs6hEKOlWKgbmZe8OscjqO+l7wTEFMmiFRu0cLBRtWbc9nR2jjPtPkd5k
QfVq/jKsJdd3WnKxrKxB5fjpamYKlEQnDpiVRfJiMY3J/Y2DoQ6PW37e7qUeYYv6EXvnDBpCJu6U
S+BOKaWVKPs00JwqnO2mrDthg3SgQTPGzidJm6VupxudiLnZpJnxBDOhIoAaZrveVd+VKuT5j2wY
rsD5eduHi4aTvB3dhtq1PW5dMaoQqURYvRNyCClOHcYyzDVgp7cYHmd6lEECM0ESb34o55zpqRm8
u3tqHO4ZiGRzC5bpLvmOeLwhWUu8DYrNN3HpAPNhdeRJzQrwcoWRDVq57QnRu4Au854h3rTlzQX3
cVFVI17UG2n4MlQSF+KLhvoPrRoHIS54AUm9UoXM3S1FLZ4aA+T7niKgFzB8AJcLVjveGhKOzUtu
13jrxQHkgNHBCRbrGOEnRF6J8z0OQ21p1/YhNDxN4ticvrpjFN6FkZ0s3Q7sYGuiZZA0aqb9hSty
Hv1tZLr79YPhVJX94r/KCSXzOFPUz53+adH+WJKh4zdJC7ES1k0hjvP8YOomP2Dl8eO+zaqqVYL6
tr+R4n5T9gFF155oaB5DGJL5KeNK3agzHK1EKQ6AOuFEf4Zp2bug4J/0hLdnRDIaWJl2VIZ5qYih
bTBK6BTpeKwNaErklCIRhmJVZc89xdtfAmNb4noHADLJvz6iWsFX9SExko5zgpH6qzle9/IMorjg
sySK5UOkv/fwrxYj4mb0DEoYlDfKQTJOCbEEzp5uJRUmskZGCjOIg1zj8/QvAG6bs/vMLaXX1vkT
24prIq7vivs4Y6eNbIVx7bpCJ4Z86lQ02yzm9PYMj4YmvR5HuQ9TviLnLFwozDRePpo7zpraaNXx
T/17KG6OF9xtOQpIkrpuGqpDCkaxYFQ9s0D/6pzeqruhAeRfKOT8ww777EvdtO1X42WHj7N5dLmr
umSlMQTwSE8jnDMlHQvbWKG3APA4KcO9Bi0zatYSWeHiSdpUj/SIPYO/9HrKY38+YtQO4jST+L3X
6JsyiCfLrEk7LzCmIw6RayU1UwO6WIVcF4AI5S8fH5dHNqyZoALNZQ5114ASqflDcDfNJX0YGn1M
bR8yYfK/9czLBSowEP0QnE5LKjL4KOaiT1G47K2LhrC84XXx/McmZAszkTjiOp7Mwg9I7iRoc1BY
Kfdciu9BeoGu/sz0FCJFjeLep2Zw0TzRm+IY/TUjYARamj2u+nJu32SW9+0pCSxgLHyRSNcJWuZt
1Bym3rmfJ9/36hBSmAtwUA6OVVWKmRAj3mm3uuedZlv7swK1Xfu0e18tkWrekXLrRF80aas7o0fb
MthOMC44Bq7iE+kc6HiwtV8X04qq9LEhDt+hrGufPu+jJTMV4jD1g/nsseEhAoHGurxFRLwMoCdt
WrH6XFmLpA2+B17QQe4upOaGkmuoaDg0MqBhm75HVlkoGjclD/Ix9NvN6hvcVuQTid6/ZF8YfQUH
rCu9hp02CTZm4byq1+BJG+lngQWrgiVkFUad9rEQFenelwus0K3d02ZqUGjIObfPPH7z2bvTi0da
hQrEuq3+dvTvWjvuxd7Z1/bxSSg+vn1gyeptlDm77eFYugqJvUA/0UyYwM9ycEmwDPh2QD51HhAj
AV47P6qzfV+q0msIqZIl7qjlwa/amRfqi0esn1r+FWDvZUJTFuEOHXl4Up9n2mN06STTav6eB8XH
PXlDedNscIPn95+sMXvhCcWracp2/3WdxDNq1TmNdEXjTLK4ORE3ZbnLQAxHA5A01GFAYn9bHK9O
vcglzpLUMHMpZ/feuNej4w+Gb11d1eSSmMnkIkZzVpSBOCVaaX6w+Xr/eijuf0dMF66/75ZSuCiJ
dtJk2XXdV5jBAGLrNByhxxh39Z9FhZ/BgByiOphIL018QdY2w40JRdCNeUU1z629IYGE4rtAacKY
VUZ/3rH9QhcPdC/YuhCqq5ZecHQWSOgtM2J3c4JpUeILsce+7DqHdLKaCRsE6n1/HSL7PercoZ7I
ApNjQ7KPQQpAeUAc98RF3zbnIQtuyodkPP3rl1vxrkBTE5sJ0m1v8maofe2C8GY3McGBUmff38hz
P16PiRakT7TSud0/5BFO+b+fBjmJaaMfzFAB+67fuFL1UIz/zkNE/N/Z0No7WHG3kKvhCL+IQSHQ
nM85d/zTBeSI0CDuG8SRBOjqwIeOHleka8EzRzRh/ELiJe1xalwEkY67LGMm9f6liCo8mbNWAlrS
F0FnNtRQRkhsgl53dX5Uxgw9bQ/2eXDQV9Fn9Yyp7hw2Kgpnsf8oHobaLvmcpAi8BPFHAjIyiyfU
E242tQrpMZv42rv1qcmxaaJ6Bsy+QnYUEeiR2b0Nc3l1GhULC4cy5mpV3w/SofO8Tct+kMHJ/sxw
9O1U54JOat48qVlpdPeJ1SXUJSI3vIPGXSiGCzZoDwkquSmzBOCaZ6R/2J8L0Q3Cuppxa22uVwa9
V7+DQjIPy5A/PUCqUzfoEmAnTZNHoW82HzU+jiqyQF8xv1OvcP8qWDWIbtdojhhVRaqpaOqZcd3P
GBQCKSbhniMsV+kEfoJugVcmKHGdGfKsbFMNkC4ejTWjDmIDxLsJPVFJyKodN8bzRZP4g69zRK+g
wfSrNemhFi433t49TEQWMoCqW9G1v3MaxKafHYRgnrgpOTS19TgwpBhVP+HWuRvwXZej87evLyy8
HK8pCvvumzGFeCNQsaiNNI/R7m9TYwKibYuPt0b3Nj4/2Kl57BAedvJ8vh8NWZGbCmrY/BHA5kNp
P7jDVmrxszTXtDX92+0SocmvTw1qzcMtKptELNAf22VcH5viSFzWiPGxcxU7YDu60Z3KeYNrlyod
lOizDPnNhtd9mk2El/e0Y4ugMaXCa0hMRK5txgo4FV3JJ9eivAhshJ39auJHqENN/yPkFSkMmu5H
0e20uspksLIauiBH1o1PNKXmwYRLSbthgVH+4Xb9j42Hi8cotVJChABk11axIabDv8axrtPUYaez
oZDXDiWqQ7GstG6/EzsC/A3UjlZQ7BYjyoywfvB7xAxII+UDcwZss/G3G9TyAmdWVCL/S9/Yzct8
UG6z9CANOmPf5fntA3lxHDMlVb34afuEfch4ECIfV7IWhSrYtUNlRTGU1zBIYNdAp8yfrmszjrHZ
6xzhwpTr7gGp6+YoGyHfb1a8T5GmkQWHSVCX+YWHP1IwLcUiBQpXNmZOr6evx4nPQrvaOuCJtWyo
SyB6kkH+0OKB6UQkBanCdCuQnxHCG/ARtIVDvFAzdrMonduGDV5kPRZrix9cNoEN36BxHilX3B2X
0e1x2AxSyoJ1kQFSo6StE7KofxHcuQi/m/l8/6Van/dHEds2onHLBTwO3ZrXs5hG/TTNFZCLQhwF
14PRsP1IUHX/eqHFiQc0jkuR+cjdu0jwI7ThnPi5QjSBKGU/ukjnirT0fa85JODSUnCXzH+/uXnE
iwhUfIzslLMKW3f3zIxfI0KdLonIzW/v4d27Ltjzob9XRgyz5ntMp+r+xhFrFlLtjoDY7/fDfbbB
jQx9BEb75KQN7KTYo0k2YQ3cRo6WCfRhwTFosa2BKu0UcUh4FCTFfu210ecck5rxNzVSrUoPKRKB
Iw0SKyF8+qE0NPB9jXGct7cQDeOQzURfl8fBL509yttbZ/avtcWop9cBgOY55L1ksY4W+WkLhk3b
VvjpBZwc4LkG0OgkTbxjt4YCnBXxwrvY7n4l3X5Fu6nj+DcdXuevgDxf5/OBJ9Paf97iKdGHjXwB
BAH5XAgr7rhIdenRgzbj2o8pCjRlHxvyuWYZ8vZCrHmryvxSyKfChiVVEsieYc+O/t6kCtG2Q2BG
tq3nK7BBjJbSAXSjRWzDjkJzd0y9ASeXm9MBa7BcyGGRZfKENE4/njwpbpgw71j8/MH5RL/sQfYk
wESB72bnkW7ZQbJQcqOfEhNtPNfFHwCgU4wDMGS3+4A5GU1Y5wMacETYOQJdLmZlP6GsyrrB0Gwd
7FiyEmOYIRVyhhmur3dxwboresDtbYvwH9xelfGS55/oIL5cgxT8JivY5P7HLelTkx1yUkX8NCAE
5QQ/itxmZ9bEUgo7FSwpjGKSGchumXNURVSrA+KAoTiuc8Xho5jvvTcMDsv9KEtIqRb4OEgWucLs
c22EvdZteDFhLSC53s+2u8/mfJI+5yroVhz/8suZaPwuC1J0f4jnGWROu5G5obw2HmthPWuxVKZP
eqpmH3F65cWlIRx3Wrh0TMegyEBM8khtYn9qRen7zX2ptqodbjGIIGuQ1PxRN2WmGEPZqxtHcBIY
5lmrCSJq9VgIUdWeVWAUpbyK5zuDvSRGJRHObaSL7u7GTAti4NE5/WgUFUpJTQMq7A90Z9asTalU
NXfrhlcjrDB1/hTanqD4tChVWBMKCPftcr+EBOZPItBjuuJpiqoSXYzloFtdpQllWxJOxbFCKpMm
acmdYIK8ZNaaLfSSnYDS73H0vo77mKLsk0FsbUfQYHcq2SHXlPejic4LWprv0nipJjdttwwGmf3d
szi69EAasq8OM0akvHJPCYBo9qdZkNfa53oHgjOZlklubnu/Ac/ddDoPbGWn22CCYDE2TNpF5oP1
3u018SPHgNBUIHou7kcdMAVRA2HZugJECI2PpdhQzYsFFOhiQkMUitnJTPiM6SGo6NGpkggMj7tM
rdC0tnvGQMG1u//qcavWeT5HCQj32uPLoYjH60OXucd05T5YzOc6AgfJi1kCErNA1UzuEn4I4dD0
KPQ9W67XYzY5UD/+xbjjWrR7GsY4KioFC4DLcQMCooqQ8bOMeWzZbtHOmTxJaiDfnr8/CKumXASJ
jnxIUZtrQP5eMhDWd0I0xmg6FW0Wiv6uL5MIBIwFZOR1kcgCJ9CSK30j8GMTU8qTNaxd/cr5A9Oi
vw4fgWVmxdzIdyV3QGrpN4SAof4tkohFw5RuE2u3ekgnuSfsD+zPOSGRzqH2XXmKp+qd8a8lZv8s
Kz5gHmrjRdR7QjRW4cXo50fILJDDR7kb+dxXXZTAiaCNIloec06sxOLCVAMIxM1/z8Ad7YwnmFMP
qu0ntMKJMy4ISLahRx7DdvTh6MVndL6M1hqf/qR3UzM/fsxVijktNDNKGHuRKZVjCRZEigRE2ByH
uxdTZOKCga6ewfwb8AZ1NYC3b5NSrGJkHl3uCW01Vo7KM1UKGg/xUUFF5VShy88Xyz6MExE009jm
jaIYzU6KLU39XUtEE+yLaBKmOPHMYTooJOegeomViBHrHT1hN1xs5ks8lI/P713HDhN1np6MQJHP
q7Gw86gsp8IiQ50o7yzKJ8uLMMfvGtCVD5oqSHIw9ZYLX9/EgdRFQAyZTePGFNSgHfRxJXLGhgU3
eETXg1pUsuts3gV0/PeVEK0AeNKOrLyW1TTT7nZRRDyJKiZzGI/Dh7HKzvgWNZZrmGqUUEmJ1Xzq
Oc5YbBDAFwXjP4FoZdWlazgxSV9GPQ8keiHcPBX4falhWPWXNPk/xGhwec/q1loP54xh+jUCa1x6
JhiU7BNUM9LAXViZ6PVF1ymFbDjFRCEeLyIEYJhgkyRThgY9ZWDcQdDLKdr2IfjavX8cela7bqHH
iVdz9T4bRUIbKL8NcbfgQfiZAkkL3WshPinpYY3d6ZCupQS/JGqU1ho5tlrDxXP6uHS1ZhkW3WHJ
6aZz1KtH/rveJ1L9KFLuZJQXo0Rkco3LiyOjnkpTaIqn5oji77uXqDIBu+8QXOHRxLDxSfkzujC9
Bi0KgzArxBHYmse08xm6RXPwcZ2lR5rNGPNzVzbSTBCHq/II1HkTLMATVMMaCf0mE/h+QPwajZmA
/gdDx7Y6X8QBw6j3xtbIOr+zEmeNUr03tUixbeDfqzO6jiB+36D0atre+t+lqWwKwscC+kahT+Sm
1y24I0yGZDsVaXq9aLTvMbGUUIjpYy2HZq2A/KYxh8DSwFY82lyLHR0pU65LeXrfwafi6KboeXX5
2awAZuMFLW7952cEhyUrjbLfRpgSCEY48kZpw9cjDjXFF/YYnYwIGc5f+B+3bA8I88RuA+DZ7hnQ
GJt4GHPCU0LzEvmivkFWBa4q+FCQ2oSRTIO+o5B6DrOv9hUb7wo8mJbD5nkC45MA3J+NTNhhUS8G
wzufGP1um26OUrpKl6kljjMcpXki8wFDE+zcKhUqZdJQNMn5gZOYjwEi7MGuHyvxkFEDRBfeljLB
jT7XRufYcA7bGyUFazjVorvDLFpfKBB4LuVV+PoGv4AyGOMxHrK1JjYouayrxt5qhiniHS7zTgOB
YtzVN3xloThU0pmonGocFZuXYQNbh2xGcUZUAa/nTYxcYZ79eYVgfKV2ItGjXrbXNZPfBkjnOkku
+alDXZgX64wvRDbdhxvcKU8AJ3VZf94PHp75M2/1rZ8mDQ4Ri+kY8oUx3VtOypPvZ3uemC7vr+D1
sDyqREbcxRaM53pazgCRJcxGgxGNlCQ9WjBEX3IkkPcQWMKuCW3JkFLV7FUvUXCqUlFcBy6llllT
54jVdrfuOulC8IMOwcalEeFnra4sFcP/s9R0VhPFkhIUdMF5X1CD2y6aRLBCGZEL49OGfw3GpVBj
b79hCarMJG37r3kVKwiIsuofYCm1l/c1o92ZDbg57qxvQoJbsYM1f3zxRBDoHIZp+SNSz6W47ffR
GZMoAn0co2DEm1TfKYilSdrOXWhJXEpFhY/EW+gr/eO9NBe0fnteQye0HJS+oUCFaCabh4irsrwp
GjnXi54mbiYukf+whN8vvfnRuP2qxQfvVoiWhUh58VcmaTa037x9ygaVkTyXlf0htFo87dtkG89s
xfNEkYJykfRjA3iaR0Hkj4oS2iseaFdBvbFvPO1bCo8FfdUJWQggAw9ggcs7gU5Wmq+e17ZJunoh
axoLUZORPy6b7Pr6cfYwowTJICC6O6GzFcUbaCKmZJHp2nvFDCCSd6jagt96TI6BNtIjG1nLhqb8
/Ex6cIBH5yConTF9/01+slUaQt6yDw0m2ME0T6D86xyJaBdrKRiB+GNlJ2I9IU2z6nfrfGthDHQk
85Rvm+O19mbkbvkHsryOBj9caKwoSqnoA24SEv7ICb70yYp0W2YMQBFyaeUJpQ7rjsb2xr5ORn3m
X/dug1ahI+PuYHpwmANFYLpLikgaGAsxvyAh5ulhPXHlSf+45uJUT/2ShsLXQ4DINjt+s7Dl9j/6
8/Xqwi6rs4m7kjzgvIG412EdzAyn0vs5dwI7Fat199O9IiDEH7iGe6t2uRbhOOobZ32LaNHH7wCI
qmdX3TQuA1RXZBFgNvWLzCV1Jz+fTp1/7mYf9MG/rQLRwEWE+tfTVr4I5rY44P+FsE4iGXMJMenH
dsaelMcmcWntY7Bd/1skcqJb4qBG+ZG1oti0IkVVec+stseNQ6IjR4Vd9+eEI+anZspNOv6sT6IW
rAi+0MbQF2oE64ALM02QWrrrIc0qV92W9isgubYr6rdZZTyf1s4hdxIZyxB6Cx7HXylzIQSQzdR5
d734ReLcJNAVP5JWEDBMyI7O4Bezhjhcj2qgpCRpjtACQg39yUTh0RpAexsv7oWnadjI7W8kV023
fQrsqUkzc/6PcaEUVRSBmJ8NAAwiDcs+IYYq7w+TyVtzMfMcM4S5D3G8eH/qlgxa6zEC+LIjenJf
G62LyGZgvScAPBqSxYKnMubCjYLEocurbtWgOQaUwImejArVnvuoItHLAE9KidbbdLKde5qYUlMF
BHkOvc9GQzyjsfOOp1dTrwkBrpEbtUpOoHwDtgdJ1vx1h2jdDrDtO2y0qghFuJGMDTvpdUaBmah2
yxYJgzROOJUxK3p79SEmFunL/HwWJHTBbTXJFmK2TtTD680FW+/mUOy82P+mD+KuAKv7X0Kd0F1B
hvfV1XPhazE46UjvW5ZbuELeXq5wsig5i//PJWNUUHZ/tW2Hcs8QMSnGkZkbS5QhHYx3n9Ujvttq
VkAMGtuqjcJqZdjfErFs5W8wjQ/ntqMvf8Yxr3WaSwe13TEtMLFclvP2vF1qmuK6JoIxEQxdVtmN
hg6Vt17OY9mryrVVEbm3PzmsJNCQ+G1cOHtGjVAi6DNJ2EsDpEXZi7m3W9faqYbdqAgynnKarpfx
YtNmbixdbyfBy75jiKKB44IqcosXaS6Ethi4oZF0Ftd49iwy1ncWk5XvPUz9LtU2K9lSjyr+5HGc
bolMp91u94VbfkCM1TnRaF/f1yboqMemXd/rqcCsUmKCgNCC7jYVIKws3AMebkp/3yOjIAVLs8VI
W1TXERKJJgRbZmIjnu6i9/JSvdue05Pb3Qci3zT1nSK/7Rscmtu/LjXSZ0u7M4SakVaTSzRgrOAz
peWElOWBG953e4i8hwD1m6hScVY7sjhl4b0P7Gtj5zbg5O/vnlcw2TGjJOVwrgVgksVG3OOeKAdm
2N9uzvYALsbMj7T77KXFxSXWXL/i+FwdcXTZgLIOPStLmjom0dZ84/enFPS/JmPO4va+6dD5ddJ6
1jxQ0vQ3BlVhLxTL6k7dPHDQWjIfRHJPuVWnp+SDRltcMzJDKwJjeazxIYYtN8qCnd7CeP+zeVSW
1NocA3V5yfX7qEOsEz/enyhbGFu7LBYAH8Zr72XDC4uIPL8U6Wv09rNFLQROdn3rdas38D6b5Q+X
Wt7y8uxOXQ7f1jxVgTtRiFhSZfULHyM0+HNsoTN/a6BTX7ON8CqGq2aur8uq47vKWjX8iow2ndgK
mBGVlKMbjo9aP+oWV0XalvXoPjx+0gciWgCYq3pMF7qUVs8RXRawsQCbc3nToW2qpgn1nQHGJ6ba
4LwTEdCrXRKlzmw8HVM9mWdK/yXPt8Dp/8JugTRpPorgnWASQjIutBvuBlpy7nIfhDwkVqvkiH+w
pXW14lHSetb7xtzOgsHV8Rxa9uipy0WkHIqpe+613cRLouOCKvLjZJbIj8JM5OdxtKdJGHVfy5yR
KduFPDtuyjVh50BL4tGAEp62n/pfOI5iG9mTTaFHFmU0s3lypKMsI/pjI6oLOvwDNHX52su5JMWm
ky8BdEooqJ4AQFOhsj7XZwnrV3yMrPWZaw5PZQpLYO38OMmGU8QN6DTTktSfqCoS2XxGcT4lMB9W
oCvgyhatOKWUh6eP7Wh8X2JkteHmdqObyqRXi1AOIOan7wL5udqftFfbMYrrmRJ/yq5e8krm16Sz
AUF5TqY375f6/wYSnr2E6JNkNUHVgFQx6AADeGGg+2lGjRzWYFyf1d5aru0vAZZ+Mdyir5QAW3ZL
F45Ay4Nn2K4e8Fe78c47c8v6/PhQgO3aMbCqjHPpua6QNlS9+posvHWNaauOhPpEPRYBRawm76fU
0OxKlNOVpFDdt59ctrwvNXh3rIYq5AdjkMbJpPppkno2U7ZfDF0va9XFd7qFOstTYGPNo4XYDTzu
C1YvCZiJF8oovq+hleZ2JyHQY0ST01qxeTyKHWUj/cwqB5VyY/BeXct8pUMvZg/u2tYf6VjjgxDb
P9oKTCUlGxxF+bWSNfYsCGxOaul5nIt+8KJX5aVqMPUZ/TTttDHDEJKOXh3mNHmVfNzyYHw00UVr
3HVdKqwLYq7F4La3QxQUaHwQXY92luQaw2qDwIWub/xLql/rhWk8/f9/l0bMzF6Yfxa+p9v1nbkw
mHLB4GKr5XHWT0V8VkXrLfJdG0iHOqNbtchEoygVnHV28QHS0FIVPaKdHRq2M/2Ni7X5HTV2zV0+
ZatL4OJ0y+32e70y3ecipWyGZwMXVgwQnKax5cG7ELtMLuFOny5MMlin3rmBmrufzDcacc0jZsmw
86BCP4EU+A5mXAgudsvvbdTpqJH2b4u6DRkzwyRDZdJCzrEb6PGc5Qu6Z1MjVVIfOqMGKhZgv0aD
Cmiwg+f51vPdinLACiFUaXPwzO7CqXm8eJEOt751MiKirVfmx3gdO14nk7C14G8C888jyhddDeiV
08tEhthx6bGyTZD4NYVbPPeiV+Bu//epJIdivCS+MNCdOmlAxklmxpiADzqZO96cmwf5eLMD8iZn
d0ubYp8KMlV+OcKVoRkloyCCswWZAg4Pnnx5evGByIsMn5gBxyiw2W5v0bfStH35kYPzaX9XxxeD
+4l8cZ8+lPW4YBcrmzqgqltc94Hype1xhSqBIJQK0rqAPJ6qyRU82Otlu+tuXLrjrTm+Uf8Tc3fm
P/QcmdU93iu+V05ESLdyhBjcMhDEY9OFWdciOIiLXNUBSaJAIsqFbi0DR+FpKp0vXmG76SpTZeDT
aV1IwU6m66BzhTNZla4b7Cg/kPOaPqGwQkEXxfEkrmMjbNwyTtdsZXxEnMxTrxE/Efa0Faouw8MT
Ya5reVs7MH4N0QhFlv4IqnJp8i3cYFECiC2/AcgG5i+mzGrNW83j+jlPTkG5/7chsZC8taAEapRs
tBCJVl/OxQtegGlBVkX0Ays8+imNV2QJ7AI/aSzUNS/RHi4LQfmIek5aUlxinqKINjHSXScwirWR
npnYekPO6Yuvm/75t+tUNHBahWgIq3Zbsi8hRcXDOKuGPTWu3QU0QuyYW9cuzqZGIJB36dBk9y2L
f8eLyOoEfu3Dwpx15DPtpuw22LkLUTpSeRIbqkf6UAT7rcKcANOkf2+2LCewDJNOtPZZ02VheQg9
FqP8dxEo+RQsx1SiIO/IwvkG1U8UGXFwbFJxKJa2TP7L2VKWW0bYrp3NKgm7strfPZ2HkkuyCO16
6XeA5zLIGz74JLFQOpkDgxY+tbRRDttTPXzLbOLW7lV+36xez5QW0zGg4yscvNACAnzUDhJG4vrH
SnXrgoWNmSFwkU615YpTwVy+854eqFeKXj+QEvGR+n8zCQZraL/zTc+inCAA/xm7bnNiUscOmQDF
+1lDnaZFqMuAvwfNtVcGRHNOcSIftWBsyD4T3g3xjnG4ZNNTnYlWD2zvYWY+hZSdI1L7z2qU8XEL
eUfEc48Dr9dVdToouUGEA87gV7mcWXQyHE3rHvQrfutfKTixSiIBUkayN0jSNrb82tntxV7R3v4M
aA+Zp/bmNEk6UnrjWZ/4z83cGJwwICc6vRujRHVYKxlWK6J/k5wvnRHsVNrCdWl0+x7M0gRvrzy3
LF/rcFEG+r6P/bNJRq7JT1nkpkeRNSEAS+ZNho/GeP2UpeerRZ+Z1X7B4CbvbgiJ6YdDi+MKluoh
yhl6YL5ZaVRTeSEprllm1/LfiASO9t/D3ax7mIDBrRKVfk2mVj9EOcoimXoRO0NkGez45DAbzEuE
UAs2Cw5ewdm8y2aa7zMoSrWqhoxQ4iQD0bHihcZpvkl1KaCMwHlMx9VXGkiXZfF7x5SQZlaVpkog
C/CWduzh/y0Pc4PhpdL4NsHGhg+rJo9n0tYDvYN0iLnEQ47AveGqU0ogwyouw+JQx/BZnruHCCMK
/OfLYMTE1PhT5H9dgWuq6Pmp5VCezwpCDihE2A9+FAtzktJgRiEE3RMu6OYG/Drr5IllEV1MxiNH
VMWxgE973V34oDKKiiWTCIRn5JjIaRlUoUOMc2mUcc8+nT8rMsvP2stLNMgtombbHVVYfdMbHY6F
fWai1Bqt90JGste6PoKnUvyLas7G9yQTXKT/xr0HI0UHa6TTMQdDZXBVONC+Dyd2teZZvJD+GVao
o8FpTEYeLkQzS2tKIYgdw0D8jWoWlBpj3//Ra7biZ0lyojEaNrGt9hzYtlY6HBoM8A6bwfcZieAR
k083R+GOxPwxhoi/aPeGkoVqdkT0VChMJsk7AXvrx1fjVop9kur8WD40Pp/SHz3zxiGMXNlWDDHn
ZW+BJL5/wKMyJdxcz11y0TSbnK5wmmji0sH3EX8VWuyzOK9xlIpaHYh1bSuYD30dsrulDYzCzKwN
GAynG9xtTymc1IIbn+ibjQHB+i1OGyu6VnNVBRKHb469DDwEIEAiP0KAnDwilUeiW49dzQd+8p/4
1zYR6L12Gw/5bpnNILzhugZlEblgwJ5YQMKvDMpWwi2y5wF/XRBCZqJnaJyzgsHECoKxmhLpruBk
4PGv2gOrt8pO2oYF4ah3pjoHNjKO5TB44q4cArtl6dNytBh4Gl8/MbvoFinf3qtsBgCHcI3RK1lT
eGFx7u+nW4H9ZnkhJziB8lKitc1LMxG/q7Pe8/wLJyhJPlKqpZe6Qo4H3dtMDwh61yFmO5ZhDUOm
eAq91QY89XOBkcBP0VqjZ9D11NzsUE7kOzih3BWackf6BL7DEjuRXYj8aTXZIINYPaK3L6JlPcqm
CtzSlAoEnevOO3SD2Ytk6zJjHOCxPNHkd67Kx6pJtLkk1KGMNN+b+tqK6IbGk8I7yoVV4xag+Vyv
PWO2wT+rWaoZAq2UmVeUVVgLJIZeFSAyjsXpQQkjb6utawUlsc6cruwKUCE5LadALxBeuEPUmoSs
fTksbt/Q+M8bk3WsMnR4jpjJQUAmUgwmoBChe12+scow/xK2qDm9+UNutfydcLqNsiA1U65kqAeK
VAsgWRYPJUhuDikuYyeCCYoXZ8JfgAg/fQi17Cjyqqld5vURM+zyJNEr7Gx4PrhNndxa/U9TrOaa
24AqVDoKOYdvFV51B6/o7Qrd/FLSj5tB/KaxkId7IF1v+T2MV2Tn8yob8Xnd8b/SBQ64s6+wBRvD
9iEORBub9WJDzmJyCCQjF9oNTWMqioKs+s7rHBJ2pA5lT8VBCXxS9YzjQyZpmTc3VkRCzvjn75Gr
YAfXjF09qsiFmE1pqTFj9aLeXGn6f9i+hdyXnFB6VfNRI1NH1IGpGl68B/A6i0VW/EIwWiT6XF8e
jWzwsMpYwyGxUAv6BNYAQzbUXfFEDxCfkKPYhgi5Sa7eXl7+HrWx/fCSZJbDlYk6zDnf1fs1XFK0
4WuZk0/vf2aPK8cY4mjgvcOWxWm87aTwIKJuiEr/BlsNqAoNzR+M5tG2S4Ioh6PH8KK/THhU1//8
tyzarqQYW8VrKfJcGzKadvlt3znWSzYivt7bM/RQN2VMn/Q9shyIpRt53n5R6WHSZ947ryQTFx2x
0pwQZlI0IbuAFcC5tf29Tfow+3sbjosPKJhse886bIF/JhIKzwetsf6w0BfFdaIbKKgse3SgEJPy
qSVJ8DBJgO4XsqFk1jYkNQJtFQBz6iNzJtPn1wPS/mN4+8v+wYVU+QaqvNG4z7kMBoaD2DZufDXQ
rw7qdbCVLgwEk5kdgPAmmpr8faTB95QCafqbHPZtTX3BmoAFGrBqXNTK8EQAffVzv+WO0pazxMk0
RL0QOxi+uS77q0ScBOVgMFJjgR29hbsbUUG8tWrA8IJAJIu1bAhJLdmiJkClzE44qMNKKfiMTBi+
TeWLOO62IwqWdp2X5g/D94eVhAC+5IjYV4l4E3nFK+vdM34nAPR8D6wfrMlb16bqrHS895Cqej/o
WLPQxqXOMnn8u9+m5wYOdg2ZKwUjQCvSGha7jkB3EqG69IEF8tttuP0cqt6pw2W9O7R+9xHxu9dO
yQH5dXUZnsJNmQ7JOoXyRsRWq8Aw7F5b+FbZ2OI8Bt0vBEsSW2Q06FCh91wIHmgmsUpBJMX8LwFo
i5bdybkStFLVkBpTxA6ac4x/5VtN5vbpO+9A8ETDkr8ag8LQ9V9PWzog2paMlDp90WIkTGEZBu5T
mXt+pNIxfsWJyM6/n2FMJL3kuOEX52+fKRkJcrjMqX8JRplQSdXauRTSt/k1JqwiGe8o24vz3Sre
UOaPSMofQedeGWBK0U/M1dbByAw1DTv9B7ZRK7J5F6XeS79rIK0Am4W1jsOZRYuhbwW4VNv51BeJ
skAdIzVGCv8PUBszMpbRhSrA2Pjie8Nh15WXg6kJBvrqPdXUSAQFcmUidfQRnTZf1umJ7vZaQTkh
8lsFMW33KpE0ZNCuPADDnX0A60TCwKChCxHneNH1QdPYpQ+jEfXNpm4t3dg+RtLen5JJ7kycWU/6
EYpGWaPRXGV7hxK+5WhUF2IEEw5Fn+nJnw3qSoH0Ne03rZXwhEtRRXP1cLShuj9TEMRBMeTtpGhi
/FSoBwPrCpd7/yUZ/YpDlbxFyxr8o/9RQn7C6cnMp6ZV+5iAHgxDlXrN8vlDdrWePPDcVAzI2Ans
bd7miItAk9y1lnljiZ6zWmzr/DOu0nq7xylRrAaeNFlrKZcP0+D+lTXkhPQajJ0lYPot54k3zT/t
ZMk6pGmSpvLBFgS+B93Xo28kDIbxz8xLN683sOcIAw0mMhNwMIqHTofuVtmqhAzMQqr7tjIt1cma
Ot5YF+m7DP0awhgHcVD765quMzEuTt+hplIyqo3/9VT6DsbhNX/h/I5hkEIyIhHcHxVhkaoeYRt+
ToR6Y0ief/abyqoka8TZqAhJ8VdlrIgyktAGWF/ZpWqGdDyrHBh+5ng2/JubFLBYajVnazMVOiyy
fnYWkY15VyAXJcrBN4rYTUSRUcin/3RzFESyuXkh1CbNkAOOzvdJd6sawnYXfDcFMYxb0sYSpo5v
g7XpZ8vQCtvq75w29GR993+Rm1dlp/s1kySJ+LMyVVRtpxI9+baQ39T7/mXnDqXgWP8oGUogtiTg
ENq39f/fWVfiTBehJ4ytWp1QGn7morWU6iBmZuYI3RJP2NTdNPTX8yK06s765dKXlHKFtIDsyS7T
kL3Th9BisgRmx+gLHyzbZ+o5JlAiM1jBsXx5PmvsmyULPb+G0jGSXRI+WcmHK9TWbMrbaROvhGA3
sYNaK81MZYJS/2TYCy13vK44pMSZQ6UwzGDfE0a67Ek4eU2B+rb0KRSZWB4wMtE+XVvPdhZEry2a
FJkLUy3EdJE8LQ4ShtzKgrDpPUuxj/p7YS4bOYj2bdqc+8X3tzMt1xHBgBzJrGcZBJ8plU8bfqe+
+4CSGTCmeolLDmbgv0OeS8aw+HzzFJbZRPIJ4Flli1oGRsk5FRGnn4S99nWimoy8yW7GWm99FwlJ
7Wh1yDLV2QdZYoWAGEiYCY1roimeR1Vhjg1+err4ej1L6do8Phi9n0Psmxvl88HCUefQlse9pAPU
1R/+qpOrVanW8wk6ZgC6eBaLuHOF/bn1YYUPCSpv5T6IFhhOpsO+OP+rr+bWIMPao/rdBlbY7Bp0
IsO2YLBvvJ/lRlNCsph2BU5gM1GVSK9CcYA4yoQyHZfXcHSrrLIg/IF2jcqeip77BNQw0SvurYE9
SwouYcqWUH0LYoJfX45tOxJj8i9uyTgyBAx530GSzUr/fq7kp+u0fcqrOP0fH4k8zonRSVMvwfZK
L8SvbDiyVk7haiX1LQ0hmNvs2f9Xag4H6b6KuawehbSuQpLfr4PwPji2C3LfwbDErAkrbpey0Xf1
xfu/UygfyXH8YGPoYzTVwtqWvhuHqHg0FStEYQSOM9z9B8MfApxUUFf8fkL4tL+FareXbwiwHHuB
xY3+l8BCz6ofTxZZDFlP6v8Ed5uhJPIB3X4QmkAr6AaT8NENMBBnPMBqP3415FM46YXYwFCtm+dR
4vquFJoOLkyWgrhH7ZHwlnHrtq51he4QAvsLA8Hwa/ytmV8BG9Pd6Mx/rGnRBMZ9wwHKZhFx8A6z
pM7eu6s/K41H98O3/gYmhAxUXBm3cygL3s+o94oz4QRC8kI2S7o8ctHpqLrRx1sxXlrAr/95Y34o
aCuc9My0R7gR44Av6nhjD+zMuCPd9pTjVaVr1zLp+h3Cm6GEQIGmDFacDGpQdYNXSGZ7gsdsLooh
zVkfZ9jj/Pl5CxU2ebIi3JpdaBooE1g2NyKs/Ue0VuCeAuEN38ff4puNWos9ZKOq3Rd2HH8jIwB9
8bwILmjB8W4xPaZ3daFUdCf21l8I7/Wr+fsHJEL7Jp197N5a/mpEP+Du2SBGa0DKh4PGekB/AOJ+
MZZwR90mr95y7LmcX5TL0/G38BlJ5eqm1MLRZ1Zan3+qVAy6XvHW28mZSD2eKdvrlXlEnQwg70c5
Ue0GSDAGNhFukMMUdsWoE9u1frDTVWwKebIViG7X3kA0uoIbESzuzpU67w01xV/jZHYYP92frXkp
OQ+jWSy/Rv+bsdvpnSWq/uwPAQMRjxhxZoWH9Sjb0dkx4V0qQIFHC9BSzX89QUGkpmnvw6utIsbZ
Uh+iIDI5VTfvJ5lq3jcrUOykdrIAggD/dHMZluP0rcVygB1dhUfCDMllXeywvlhqzFlZQM1JLomt
5Jwzw8EJ+cxy2vpAYYLaZCFCg/a4CRjQ6hnWrxyYBuo4hx0L2E12xexFRoQaFcMPOsh1m844U6p1
cobbGUKatGO8qL/oc/9k+jvGC5DGiH3vg/kQ7Ge1MQN4sBChYaLyy5TsING9qC/4nRUpGB6KjrpT
hAmwgKndDhJjNLpUcxfuv68pNvZl+mjePYQXpzSFyt5EHFxn5By0pojei0jTm4KvdeYt5xuFWmpu
IA00erYujuvP1rIUK7AaT643yGwIFc73e4F1pizfAskxoal52FhW7S4A2Ne+ub6Mg3x4i+E/8ji4
HK1PfoLpHZZqYqaXGqF71+NRqCWSa6mq2vu8UB2DNNwSKK8LqM1n5asksYQBqtDJ26SluV9lksbo
TP8YuycJYsKtCnuCxFEDrIuwXz0d1f648kQlC+aOW6wevY0uHCpVJoO+8yBnRH9fPBFciHiMLt2y
K/Id07wjFTK2Hu0Bk1PQ9eMUGpMaClvdfG6tVA+0ONcn3cKvjMdbX6uremympR0a7q3nvtnJvVX+
nidR/dj8aZP9r3rAt1bFsSX2BlBI8cAw++lj6+tRrRvMSggnfORVlRgQD9Cg56TF1oiueT1lDHFG
gkJBUnSJdBDNY566FxOF7aAI5ktSK3JlQloT2WkHHCrVo25K8C0t2pWw8QqD4RSnc0JHglnMdFNM
CgXFvFHIWVLUhKtnlHlOJ6glIHymlodhS+HZ8C6Yj/XUglhyYYKXRFuwW7csD2VCJuXvG7KGll5B
757ZVypD5jG8tnB6FBP1BGSuOGChmI0A5a7US6VI9wk6bfef+KphWAWzKPahzswyE4+h+iuwGTfA
EUYUqFw23YmANO2RWtw2pFxaM/OIxvzUA4+qgsNVAUqrXs1PMo4eIcURsqN/AZnqfto9dMN71yPl
NHkIRP3BiXr+lJocn5qeYugicSIN/Ts4dKB3u0TkXgvb2Tk8T2NS8UtiQ1HC8aZL98ml3IvPuP83
7XA4AXul/CHPQS3ha+jD99nDK/JOz4hGQBBznqfRarKkNiS+h7FiIMyR5DxtZT+ksGiMcHByMdlE
sqEsbAyAPBMHt+prfJwJzurW1kT4WZMGZTHFzY66bdIqHAC4KQyWz3BMqNSlj1P/rJoNLIp1OLD5
cOw+7i6N2j7pEjgF4RlJ56X7PLLnrjwHaUSz2HPZIKSCPgHGghdB6iVdHYFOowyIvFCPXYGQqPuU
yg645QwRVeYUhZLR+Zw0oQC0OK0VqGdLPE01fyaW3ol4Irb0ib72IbGI0pwWqoITgGGIn3GO3234
hJySgnjs9vda7lOjFhHFcrYDj24DC43Vu6LIaS/FxLCuel4NCc0qmnzNmZqo+YhCNuu8T0tFWxdW
KY0k+qUnuNDuSGl/Q+WKWXmPRnX6lh2T4+Q2wExWN/FRLuQOpuhtk3jDA2DUKXFGI3nw+C/BU7yN
wLNtzOHQBx+GrAYPNtofHHARcMM2hf+vnc91OnA5DR+PcBcCbKfcXlzWrciq1Eynq3IpNtCZgLk7
85IztVlR7a2H6jB+OFElSCU0PDrXe6rcecJ338ghjhGKfAJBALW8vCc/JBs2WuO+PsP+7bEqO8r/
/E5cRzMlNeGjMH68M73W57aZK/yvGdlKgvzOxzmDO6zfFHYFWvc78ZmveAxjcukxN3+/SFSKMRoT
Kljwc1SLkPC0TpxNqMoIYJ7qwH9uV00bDck+HdjJpKh5Bq4H/wuypQwQKSmnJCpDKIhYOXvbBue9
aveIa0Gxuc3AMaDAOdxf/dYn7rcCas374zzAYI1RLQKxTH6own10K1daM0k59yTh+KzDGwJxo0rN
j8wQ18WpOkrR5veKNUf2JbmUjq3H93EDojLm+FBeUsDkr4Vf3dKwjIt2VP0RdbmZTDaU1zwywnQi
tY6NwJAnExjO7xxQshTr/8xfpyJ4HqK1Wt6ZaNVX+zJxdGfjeRx7tRVf7B4hwK+nS7Eepm+QM1me
8EZ8sg1mSyhvPNhdWFyUwUexVNicxdyTUqCFhBTckNaqRRuFR0PFefwMLtTSz73MnkzCnvjkXTEF
B5hYhdSEmsfHpWs5ae01/qNioYmDFE3FR/+7VlhQEEh3szMiJJlNEpVzev76VEXXMecgazgsf66q
2bEEuT9RlROTAZC5vgsdnH0r9CYy5iK7h7HOMUj/L7QhP4pUpD70XTBzScS2UKRI+m/tm0fHVhR3
+MEk6qJaqbhpx/5pD4+PAv2mo74QRj750/d0P2p1la63yO0Oc2e5utYMcvOszY6GX70If0njOfQA
o5OFd3n7CkQ2hqO7Db6Yr69ZOuPoLYKCNlyybdaTg1VGQ41Txpqr9sZKn6sF+Jf4WhfAjwOXANDH
1vO/GUo020rF19kmLbi4aP3aIJyVQLWvx7z4pi51RgwFoZpRQTVOiKMJzVfmCNi2XOm0X10jIMJ2
H1W+UI8MwSIoRIxyw1e9fVnAN6dxV7IlIy19cAIhIaIgzOln4TA8Lne/mFQxlpTh13yR+DkM+pY8
VPk1xlgtYfYTrxnFva0L7Fl8p6Cv1yZLVOVdS/08T7HaiC9mLIKcfgVKsIKAMLRhSmDPcNlMyYjP
6qIqxIrujxz5SfjEY45FJf2i3KpbOum8R5qB+Souz01w0EdVntK/1iiFgcpGOlTxncb0ImF0Jk8H
8aM8vdmyLEAyYF2EtTKXPICdlErDnO5O8h35FweZIEp8dUFSZavKt+6YX4Gt/iUMO+RpCR06RDrr
rSXxs6x+kVKO+lZQX88m+N62tBWMvmorSQJnNlEN3AolKH5XLrs0nRKvMjUUtJC7LR7p5x/yxQIQ
Jzci3RrgqYH9SC+qJbxCm2yzn9+mrZVOBnCVov58GdAHhY0F1vVK4GI7mc6he7oLw3pqBqufdacc
2iYlMZsV0lDDiNIh5cjANzRmWWKTFieRhsRVL8Z7IdGMZpktX1JqjPGTy0QeQo4Ua3eobjM2dS2t
kKDE0cB+6LHASPPhPZZ303aA/EoEpbWENn2DR6vJxwaGm2zs604na29LFjPf5nvluX3insy+INbP
QBX8+Oy33MCGAN7l92v5z+fyfhB4PMB6LGRCUIlgOjChQqrwXlzEMxRtuNnew5ew2J2/W9jQelYz
fYQrSmSR/ZRLM4jm44SSWz5mReeyT0ArK2tLE71ISkHsVzveKy0u9UfX7Xe9oD4viyVuoHgbE8Fb
F7oxhgRfugCukB/nk6zy6+mvTsmH3/t36Q6EzC55GcBsFwmweg3ODwa4uDv+hKHmEHTN19pBN3ND
0TL6opLf7siKqxnYD3dyQIrQvrKFvEsxnEkbg3zPP8o9L8MnYo79FFsvF1SoXEzkiZXdIabY+m5z
rS5fa9YqQBCTFWkrw9SpGnOHmTSy39HxdfrmzI8WOTUeNuM0TB2uG+pWwdVgQP5wJxguQeHO8MJT
SY2p73+V3WKJExEvqOQDyQngEgKCjpMfG205KGhI2KH/KqI728pcoSVDKCsdqzfQt21SFT62++kR
N//3xbFDZOt46XONSyBUBQjmOGwVkmKaZV00z/Cs2CdoPHYTL+HCDWHkoY7pxfpjAWmwXn72z873
t12bM5KlqkLc4FrVUPtyVMEWQ6Eige4YW573WWo9CYEnDrxw9Jb2jPr+PmXBAG6kK3rvE2PACbVn
ayU8poLCsd2rnL14JNJKURr2AXUTpzmJ0thSgC6aQyMwHLTyR0wXK7AWU0wIc1rvn572utXCqrWV
sNqFAGg/z5kTeCAhLEduyNCX6oQSN+5LE6tXOfTfSBUvE0iZY90Q5jm0faPRHFRyRt2m+a1dBRE3
XjkujffGZnG2sRVT5eJUr2+NmEk5MBAt3wVh+eHT5N4gX4WluJJhPcXfroc5xL72gCZVxbfN400w
l2rW6vnenoA6qfxy/zamrbaFrm3ZD/7UVkb+Btqo7x8laDG1k8oRut/qxVjIAEDgzAqepHRwDZkT
/lodkP8JhWGClV5ZsRMQjV99ixv12dd5z2JmfjCz/6f/29LqaQQgGmQY1jpQ3YGSmrz5MDdFh9Ld
UnL25+Mx1qXGzplFBx2WCTCH0vOjjBy4c2qACIe7B/GiU6nOLOVFPhtyv7lRB+5rto6aqWdRKXyW
A63iYfLjpVyMMsFJmmZKbp+Q5mZiUseDf9+1JYaDcza8Z8xqMwLz2jvRNSQSGdHlCq6th0eoS0R4
wZ06XShCuM5xKZLb9tHHkem5J6MO7IkhEsul0IDtyn+j2OPckIWAt733tdtN731HNP0XG+nqRPfk
Q6XwVzzqMPQd2hgnr8PupaIBBT1aWmHgcy+ghteLzCeOa2K0MpHyg7suCvVatHJ4iGkK4JT7QVlr
xgQy9YZxZ6DDCy2W7H+fwb6/sXyKrlrRPNfKO4fWNJkE74HtR2Lp/tj0l3ehaLbGuJlaiKhhhKW0
jZ4NCdBnNk/6tQM/lK7DysBLZsYicL3UBX/YsoHrzxFCCrfCfYGdlG23fabTXBpV55WfTYafVi1s
t5cvQUAMVm6i9AbXqzBlMFzNxIrkFmQrj0+iEJmhUbDoZu4yH/YjNPHdGcNxZKqBEcl7twT+bedQ
iarooCP6WgmUZOZXm8d7j/Q/rQwjfxV5hkr26QGzkrKt6NLn0CPU9L0Op+K+sgryv97OEgLzw3rU
W44FkcdI9yhbofQ2Sdnn5adOxR6+LP8w/3Y0CzbiTkivYlCsint13yTcJxtldkD9ExHx8n3gy+ma
zs2AKwNuTeWdq5/LD5tBOFVH2ypJW9tOAsSGrWnmEfaVUqiqxvDLwdpFj+YD1PjQlT3toZ6cPm5c
QWfTqMTcm0eDcCJxqt34iDlNXlNc3LtrVaIuTdyaPLlv7gevgZq7M2jYe/W6UvyMPhx1FdUMWNrL
VoggKoppNU6csDdwm3d/2NC4+Xam+8FaHbQA4ggDQNkfxPB8qjHkbrs7ep+91Ppgmx3+jykjSpSh
xBvcY+NQ4T6AY3e59ODgWkERn74edojjY4+RZ5FG745Ll4zR5UK7Zyf5qI9bWG2ZwwCB9MvLWDyG
dvwVNJ00qRL0853txfKmHkypM4YhiWL7QUdVd+Ky2AL2qkXMnYshAblSQZRNRxnPRwIOoRVo/3Ui
dgg35MPP7MTjoCqIniwx7vG1dvdAo/NI8rpHZqzLui/e+FYMsRWN02ylkcub1gN53E3y7H4He2iv
zFXysGcFOcrA2p00f+rT20G0H5Hl2grC6k4mE/pR6oPLijtMS+KMxjUtK5453Jna5f5738i6Of6x
ML/LrQeZX6QK2jAQQa+MOyEMqDi03lCsKS3B/sUDmGJD2nuUKoorh5euLPxcu/LTNy1C8ixSu4OQ
94jlIJsgwT5Y2Lav2owTo3Z7o7+OcgukPP3aPxI6yMeLPpwtRPuq6Z2Dyk7Jkv3d0hYxsxeSoBdS
Qfi3Ky+EyPMjg0sQWLTW2uypz5bUqr+NbVQW0R/ZnLrJ7K9/RQwH6LkplwGMbfF+LgRSwgMFdKV9
6hHX5opibSrFP0IV1Z77WDiwJ5V9m6DJlaHGiaoN8N5BHP+iClW+3Blsek0bROga5PlQuQS4a0pf
15AmKIwXkpSQsW+jQ36suI0Kq+KUXChVY35+OtWjS9MxXXfe3wX0kJ814jb/BL8UwooaW2ZoPz0r
kRnl7lh2UDTv6/C1oFTSiJ4U9C+eqY4oJ0dNfppgCR9ey7hE147SO3kgTSWRQyeqs9oGAIfcDzZx
BncnSiFsOTSnP34H6JGNNxr3bkfEEiWaB289IcklO0nvMQXzfq/QpkZ7W9KHMrMVpUtrZ192ZVw4
jgSFWScXlJse8HDXaL2nCO0V3Lz944Tpb0kij3ARTfh8SPxJwzsZu4H6r79iTmyd5KFt4bjBf9DG
e4spitc3LBkQwgMjS1LwMM+hwt69NQyGcJzHhvAfEEvBAGU1r+J362+4EcS0J7FIzN2RA4Dohfma
kWe77FnDXAV6XBpPXo3oKZdn6qT8HUpXp/RAU3zDmDjSk3iWYsP7XiSBLBXsnmZVz7LYXOM+RxC7
XNaP7eJXATmtRuV01LILXpSlUGRnovg7V1MwamRPzHiKD995GjXUVsiwycuu34jc8Zh1e3JTsUlp
I02dUUVJwSR67P4Ye5jpONgF7dlkScQPg1rzAJO6ZGjYtkWK5R/yiZ6jHIu0mEh5jE/tADRLbcxe
VmyRTmtoE+oBtagdlVHibgPuRte6TjNGMruUmYJf5gq48Pqq0fOMHR7aRvjSVCNM78E1EnfEHXjK
eADMndDN3sovsCaxGkuJtOrgXbD2UyeBzPOvUl2d5kCXIBomy86BLINZ0u7InzVJGXLmiry/kDKX
IIrtWs4ox0bHX6Jt2b0hA8s70z1h4cSBU0f/JWYWDZ/AvFOA6Tdn5waq7T3ZMV+K2ouewJwId5lf
7veVsgdO2Oi9Ks5j+eBpQshzTz4vkfifkafB4v8nKrKZI/Me/xYcP6YJ0seAq73TZ1Jqop6m3NEN
5tRCj/EuvtctVYYvk0Um1ZFiKl1MDM8a1S/eO8eefQ45ow448beiMea47PbohyTr1ELUxM34lYtF
5gaB3jYV0zPcqhM71f+RtQGoQzS7pxlIYqhFsXJ8wdtYfeR0C+ufHRiiSz2ZCnSmTTm3AKeMuCrR
YzvWiMyZmDB18RmmY49C9AC5acz2KPpPykkEYyN9oXt9BUstLhc4rP/7rHznLz5ktlFHWWSbnIWZ
NCp8qvcIhu4zj1um2UCzzCaiOa5IDCTMG4ujOd5UyhI80WjWT/wsJduFQl72YWp+N5Dw7brEeYAh
hpLc3sAk/iSq5vj6VT51ji2Sq16LSCuh6o0YiGTjzNB6Qs3N8UWljUp6ann3IQpKFHkVA/GTPaly
IGhsG0CpLNI1pxMET8Gc9oF3sqQm5hY3bWHN9mGMzwUcdOMFoZ6opdPYicG1p7wLYR9mDPQ0EMX+
Jbe8mzU9/xvCGZ6IEYaNRV5F18Tp+PgYJotKindjonYDxzjx948a2DDlw51nRWVvti94vWyq8Uts
dE8H2Rp3xCxitd15XH4+ruyfSVJ7yauS7GiU5KxfhivpMwkqnogis3fbA7s0GqeULogsyCGG9HjU
9QVnjIcTCdj7G0UbAeHlULWTcQAu5K5jBKkwEFTUIZ14UjFyvYvuwL+Ftd1HJYVZzxcsOkXDIJns
0qPKr2xvu5/vbSWXCodB9Qgte8X2etcmb4UbppiwjkSfL7RdtLiMBeMPmbI9rRVax75yFktEPw0Y
XvkBPBpktmJFwYzkonJcNX2fvb1cprAdmJygwdNUHqedDKLqlZvrw8yD/1ZvPTWUT1xf/611MX/8
KObuwNN9hnKhvhCuh7JRE6zvx1CDVVdEeXPcSs8mIKkHnPz6VVBkTE4dserFHgrVUJHfq+noJyRe
nDc9yi+nQmxfsylNsOrwvIV53EVK8CwZ/ICzSOjh+z+6AjnUIun2w1qe6C8wORyfGnLjOd2FqgRt
pGtDyASc7Ifrg3LqmA9gJAcqkfcYHUsRPsF6h9EEcI022H541hORFArVu2MbLVRzqY2c51ZIU2Gl
nKhwH9TgmSYZv4joLXpsmRd1H4gc3ek+oMAUMlVFfahL9D2AYX3uCZv4dS7XJ7nxEYN9HWpU35So
CjBil6rQSUzEFt+UfVLXXFDpqfKEUSDZRuyd7x+9IPwcmlAt3pfF3KIqnT+0WZzAKSuu66+q2oFl
cFneYAAGcFdXxMvwf00dGoS52QAN62S9fBq92H++ldCwPrmr/T/cm4mGZdh7ys+OkJgx/vMY2IQ5
A6DyLfKvfMRosbQ5+JtfneG2VeTFphnCiBRmogB1gR7B7xTlLOcbet2rSxQWZtEb9jNVku0Xt+oZ
zceWjEVGHUyoPq/Q4K4gS/gYhFW3oHrJbpvsksl+kmUp650vB+aF0lsyPKNshOxd8kCNfwFwT++M
OF/NT/xYh1N8q16TZcPV/ktIb3E4vrNpN0/V4MFLY5S9LVtD3LrF32XcNjrzU2Efo6E9JDlt0Js4
m1P1Bycwoy0tM0REEBtyj70i5Kvsbk1B0XW1boKghgAA64AWVv6/qaMryxRHgq/qqpvpfYrbH+3z
VjUffkbGVwQSnqQIMxs8ztrL8oVBY2WfEqc/9JZVgtXULtQ6JV8Ozjq5VsPGwYqx+tJDE+Aok4Tv
VozjiasPUHdxtgZVkIIRzDerOuTDW+hMXUO8WdQteRt++nzA7gymwx/wtr5Brgscw6OlUaZQd/LK
kMmqP2xp/MOSQGQD93o6Kr8HfTXV+21IkKuYNuFPBTU3s4v1nw+ZJu2TXEqTQdX+PiDznaAfa3Gd
IspUx7rm77kMghXdVi+2BcsOHtfHHuJdBDik7wEFtl/mnzUei4pdhx0NX7/0ju+/VRNh8d5uHjYG
iLm8zgzAXTGmpCW+Gi/d4ACrGE//CE+rXT5U6nbiVolFXv37Ctk95MCt3mFxRCtsr9clWMLrz7Ya
e5uw4YIzCsjJJdGF/mV0Ygl3u0uJFQAPO3J5q8ks7lV9MAs2T+cFohgPnHoVm7za/H7ZwsFybC0x
iLgNigvPM830OF0KI+Yyq4maV2nwBscM1n6PP0DPdoDmxUXkmO/0F6Y6/ps0DRJ5m0wH2/Kh9eiq
8bC45WxVFV1/tGQAbwkYmMbNDMV80B5dndNYRPbKQI8//i+v9Q//mCeXDshbYLdyYo6B2Ce5u9t1
krQvslYwnIftnaNDh2pjaWb621ydTzMgCuAlfJ5wg9rVA/R5wkzKh/cUGdN+5GTH77ZTf8IwJ1ly
trTsrLpE81oKqD+hrkFa7R8pzv2GjXm9qzcerHkB6rtyAiuu0od+XfT566I7jrdQHZYEu6W4llup
QhVhVJTkHHV8P1hYeumZuyjRUF2mXTSThn1zoXB+XpQUytnvcbQH/sb4kFvJA3Yid9hLvbeKHg8O
D6FBaq7lWOQiEN6lCd5R/3H3tEscjdPbr72BDmR2+GrrgzkxwgnDZ9GE3nfUi4jcgwNpx9sMZxh1
V2H26yzHyR6fDQFNPYmgJtd557q0KupTeSNTb4Y0GMCXyc5cyQBwf1NIbGdmlkSsiGLWaFv0V17T
K1CsjnPevDS8XXdz0vVXdaGSAWc+4BpN4xJLq7k3ykXgz26AfmACH3EpS4bzGMGSRqnzBxL1jvOF
ZmJqdMTcOP8VeIRSD6cG/aeOjHuoZvW5w3Pa5YzoDY0jrd3RefqmDtx075oEsWZGCiuBBVW/LnUT
T+6gQ+b2jHxEn7y5D0fKBr80lbL0fKSau3+/ZfJ+7aa4B3mKQ4BgwvFijgA6NjbGX0V2gSaDwWJ2
cH9/5MB7UXp/A6qd94H8+ek0FKqok27XZ0QV6j54fEqsE5da+kMHwf4eOrmgMs7BhHgUib1bfwYi
BUvuT67HY2EQjXpROTjYdVVbYLxFsDgBfo7uB9Hd0T8HoBLpcZ2aosC13PxxoIEjqWL7RVoIW86p
VBBnjICQLmMZqffbtdkR08mhFpuEHa+QhqGL9WINeEDyzth/lKqH8vrG+cL/Zd4VnMMFGq72v6DX
ppFcmY6uJlsj4KkOedVBJfEQ+AFhLPFo1rgxtrJrg27zxU8cO+4QWkr0uz8ZB/A9OV2MLLV0snnV
fQyeiNk/NTyJSYbDAj6IUusaWMQcYNK8zHdY61S5g6PsNRZ+ym6rGsWc/pmNdcOmI9/YqBglry/n
OP8zRn5cy25SoD7HG8Tf/jQTTBvIq0mtEx8orqkWa8OQko2fPOf//xypSuZzbiXAQSosSmXtC/JB
aK8/NOgtKFFj/BM3Ls+1RR1iPaadAI8xgqNfuRqhRpeV/O2etLtSPLZTpWvcNYKgcYzt9UKwnR61
qmlF9SE7Uayytau2U/gIBbZ7uZZw9CqSOZxHiSOuG9NTBw8LYaE+QP4Epgvj6t8gPBW/ps0+cDDV
OhP+boLHWuE9hCqAmUb2mQ4gfHaUM+zNfzMGLlvOQvbestEG4JXKyqHV8XJ3r876ZZOroWotEqwh
b+3JXb+5KoU6b9zJ5DMQtgAmsXijgKaDo7U/tPWSbeStCIHNzDLYMKMwYvgIsR0Uhlsqn8kbz/RH
EhGx/a/kQ+/isZXCPRWku1DxcSEZ8hhjAfE8oCpf7cAUDQ2rJRj21olHI+feJ6l0mP6X/6IPmPEg
SvJqP0eRnmV5N4B1Z3+WJA9lZz0cw64nCU53dHoDemNsBS8G0m9h4Uucb3Vp74FjS2S7Fd0waTWB
uYnP1zYcCoImLuBOC7Q/HqFFEvd0CZ61/tDOZbQlvWxkb9PTBjlCh/HnSs7hPKYALCaWJuwLDEnA
msRFhpJcsIDsGDrb66pQZASql2irBqa1yPXWy7iUbh6vIrSvEAiNxxsAjB2EzE3kUw0lFkudUbc7
r0uNMQQ9aRC8ovF2+RL1S0q+NPhk9bK6y0zLHxVVuEKB6fKn2xHDma8a7715N3LZu0V5IMjH3E5L
6fH0xNtPVzU5bZtDsVISa8jhzYLcxSVqLM/CJJGdKOnseZijFnbYyDsB9FIL5TGIk51ooiupttyD
uYGApVDVoBcuwkozGLjGUoZCmfhoPnAl/dqudXPH69Qda6BOoFjNzbTT8HnDjhy8wAa/4l565iRn
KJvs1A5mAhgaK16g+KUV0lRzbtn/wspOk2jh/bAvbyCpkvwvBCa7Teb2GvzmeQAugU4NGJjCHvNp
8QttuzOqQPtJ/2mFAXKbnbiXDSN28KbINMM35tdZ9vFXRQs+XT+aqbJDL7Jnzn7ANdRwvAoCxLAM
kPlk7sJO86PQvB3NPVNhVDcigwoSMXyku9CnUg1hwHJN/Pd1fBAxhvmKslf+yI8fnM0bRLisLO0+
ul4FMwsr273XQHEHIpj9xn5xksazg8V+KNq91WNIBdTd1/3FM4b+8Qn42WdeE2ZZVMFc6z2yC1/c
xmVheOHyI/ZvJKOaz4Pc0WpbotQLf4yOcfr0GYb3yQWhkY2+mYQ1lUNBJ4aQguqba+1t7umLQLUB
L8nl6VgAhlgmvbPHi815pg3Nf2fBevt0AuuYo+ge7N6J01/DAR57oaswVoi5gawVNh4Hp5ykCg5c
YtJO3yolvUE1AHXSKIAYcSGpVQuo9HwfXp6ASVxRypsu7bZ/ScPu5ktliSjXpzu8G/InkHHkD1EE
8DV4vt/FBo68eBn5k24JfiJNJc7KaRcXmtJlvOv520lmw7qQ5QRUtctyky2Vn7vezcD2IVzIrERs
CiRbxc1rE0Xavv/e5HRHu8X/TBOzsx/6qo1/YrXSUz+Z5oRQGh7wbUkXkCpDHp4BKdii9RE6LSP3
TTy5QZDNTeUFFUMvW8LztKdJ0HaUpNCFct0WnFlL6UzdtVA1IB/bYFXtpeTF/fU/fKqVwCSgftDP
ZrJyzRWMosXPH0SM4AKcqnKYkCLPZtYKUev62YuYBq4L3eFPNFxI7FN4kVTnA/RgV1v/kgsZgAF5
4rvxhGsqrXk8jfyQu39iz38yp8UFKR+BmRcKowU3GaRjKM0Jr1W5HHkbVXBxYLieTzBaJYW6e5LN
p+zuLnTwVpSod7/PDweo3DYOMb15XHNrXXz2kq0MN+RO0DieGE7Aba/roiKMqagiRjsfn4OXIMLm
1k/UhujTqFLYW3amh//wgtOW+F4IMbeN13oWnOekbasuxlm4/2JKnP45PjT7NwUg4tl61E0nMxwW
meSE98aOryz3oO8y1nWOEPReNLqsNM0hNwYvW4Po1n7deZn+wV9ioJqbhlLaUOumtVA8ipHgFbbD
lHAWrlQmK2677Ge4AWG+IAEwBgxT6AZG3G6OUigD8NTRZoxx1MCNON/8d+i34o7HeR89Rsr8uCkP
sWdhB+SCKlNI6ldynVbe11fs6z7cmF+9oAiYZbjIlxd8a0Thq+fp7sXnruoA1WlMAJH2j2dV+mVt
9BRuno5AAfHtr8LMDSBsnh9XUoAW2z4F7K+CDrVomEXqN3rgtAbi4aDUSDUpyGK1uF9GfxoYDKrQ
wMltmEstpQOE5gDgsM9q8WU/te+PvA5TyzKno1JsKVKEBHga+WqpHs7v+u0IWOu9/rOhY2BytciQ
YqE5fDcHsZgJ4zaendjoVb5Ds1zQj059p4F81QQp8hPrLAihBvOd3av/REX0eqVZez+c4NREyhhf
skK8h4Hp2cyInwHqOz0tZzmOsdA3LiF8DNSL/oTM/k6GaYL05fgQ5EVKRgSfqLPmiKO7Qe7VQcnL
gr/jnuIauev4oA/H79MaMcqMBTfuAu73862PbSTM8SA54hk8A8njp4iB6tIce9e931g90KYUeSaY
MKIff+ePuyaF/GHMyNW16g75WxDQHrveujXM9dhJKydQ04p0V9V+VK9KnEFxzVUcvZpiie9ZGQm9
bIzF3AtrmUH8x6eglK9krucSZ4LjLXvj2LuFxNdK7SzQy/tlq4N12Tf0mgTvmXL++/88hWACSqFF
B6c1sEr+mOhz9xf4P6zG/vGrqelk1fj3dC6sf904D7R4hKqrDtngMxH1k0mOQqa/pOWWkdDP1FUj
oizUkcNqwNp8bigadGI871au8+/4Boj9E7QRZCBsQguD8s0QLvUaibs685yMhnsmCHiQQHQqd4h4
Cg438ZONEN/gM4PqLGLvRQMQdd8wT2HgMEZlcLayDNrylD1D2r8zdjhVjT5OWfB3zGWzelNMMZEi
GOXBFmlYpopRKKOuvTMdF6Abn5et73afl7G4QCgd3FxMYWY8wTmGDWCpJ6wDsy9oFzVrTyBAxqkA
oUQDdo0eotcHps/aDON75mpNRSs0SVZ55RBpjTJMbPY2U3NmfHvRgUTb/Ts3/ndRcV5BTI/3VC4c
R/OPq2zwLiZwrzNx4Eiwu42obmHKFfazV+OqYk5DTCCvGHYMHTWKLDNgSXhEwHXj5BYk9KWk7aZp
lnMaggMu8u59xDRd6DFWsz9kRMET08VbJdppzz1klZt7L1sNSgizOi//ygxowt6mtcmOfX3Bo3qG
RVrgaMaNs7aW4mGk/sbjCEsmYFrDEbmkZ5Al4iIL6i4peSTWAgPL/zTLUznWqBWjUDqNqs/WVwlj
+q3u68mXEawC5h9FG71n5V438sFbNJyFu3LrsfGnB8u8RFqHrz7s3gcZOVUv6kNV+MHvW7G9yzMq
3/Svh83i/w8m21WUXxNV8QIgMYb0gh8FtEkUzVLEJ01Lk5liUbHzYoxOBZpcu/ahNqBfkA3sIMCZ
Uiga26T9vwNBkB7LVdeJlr0QDXS5hc1dCmx+KkR+/clYNCH5ygskCEvdr0p0VlGJhyt1LR/E+PUP
ecKj2mGmj4ZdoQgeW62erB//io9UKZZvBpE6NlOUMWtjtBSaxHn+YCSMYmEa2cMADruQF/lG3+eu
pwPShJt7YB3rHkzvlKUOuvijmQad6sTvJa+dTiYubGq3C2Oanq29ccH/NkNGBuDXxuy5cVdwcyV5
Emeie0doSJMbUZKGhiTx/BUswoh1XeNQXkpLtP3cgh3O9Rbq7B+RD3vu8DqE4DicNgZzK990IVyy
//vLBr6WoCldrd8Z1KQUeI2qeojN6guMN0pHMQn3o716pgT+JlOgZK8vH9DPoOHva+nneAnL9hkI
WWqMSvyCDyDV9SmUz3At7p9B9BJzSsrqtVLhyPouvjpd9wbsG56+EDYg/Ojyqy5E9QEV5Nl2arl5
nd7GkTo2R2Dt6N5BNXyQGHtUirbxry5WyAXPV3TPOKi/03bXG8C8j+OeG3r3tLqpsukMl7fo3YPb
CU6+ewvMUWeUpFi4Gb3GJY7y0V1KGExVw8fheuTcZNpR+QOF6YXmoI2K+CK1GTu8DOhU/mvXSNzG
7qrI7fnK7OawMKqOr1kHmjOYyEABi40pIK//DU0xp/0/OSSIY7WYmNUPk048b3s1x3/dYlkJVg0u
Sk3JIOu2fGRqpgvUMURgvrpe5y/x/nZw/uFczGll+Y5mKhENWS2SyFmtsRSfMAyW9Ts7fbRbffW2
4T9lkXCaCYCq4qsSwMbdpM2GAgNb2zgpwkNTuIvijRRMLC66d53AbzOAm87nhG7bdgUCObF7F5+a
xKsdQhqHpiUlUPjTpouI9bPNslP1b1ynQp3CSFHWZVvrsrceQhTjOrPscmVvwbkTafJi4D4RjYnp
dU0yHfeu4lbfgrLnxSYeOJqcGHOyNsefgrj7QW6Cnrfyd15qMqgri5A666uUlaINIM2qMGuEvUWB
uAMkI9ggO2pQt8XuxduicpoWeMtJ9kBXC7uG24GQnOOwI2Mva9ahzEC09t1aLiXKR34uEJrGJKHc
6BXUm2sKiiyrpakVubjTwHks468Uqxn6ZHUkst6L8jw1RIkZ/msA8jOCR9Od49CmEvCm5eqdm9kK
gvNmvkQIjstsxovOXkrcm2LoBlfpDLwBFYH7wFFZ8r4q6g+uLKioUuq6aF2bEfcgWrqwoL1DQTcM
SXRiWNexz1FoMzohT3VxZN6m6ZEXTxLPMj/99NHzbfimRZ+p3aVLeTJSROASXkP0uTnisfwYWxKK
sGqZrfJGSh4TMWHggchXvAIdTx76/CNjN+LIhHgNyzqEZ+wIokNi8jYe5lz82/E5BWvNqt3tdRVy
dGDLNHuKHzBFqOa5rCq3xxHXdis/fxWdV3QNNtJJUJFNmOCrKJieng9pIU7xLHloUCCPOQMDBdPH
r4jzu/ugd1+Z7ilfIgnMJSZYgw0EAny5f7+aJ/EB1fITJg8/rbtwPSbLgBjlWsKrKfM0fKw6Z4LM
QyNiyaA0JDtvoRqCpoOvovo20TBFKaqn2UlPkMvBNZOLximXUm5KM/ZyfLhHO6BJUdGJhiVjbp8w
5WU99iZ/RjbG21KbpG5vDluvdSWnlH45xGjE1AvLVX7OvCDbSytzzH0pTbySLWvEMFzCCFz9OSv1
reR0FX7Zih+zye6olxLtVB95cFipmXLez4AfiJX7UZSjwU4WdyE2OIwSgy7hu2/EJ+T6MtYXPFk/
MhTdq+eNEZET5csv0vCSHNmo1MwCmw4eNs8yYx+k49rdrBN5di8VMttjLJe1g4DiIUJoDTNigC+k
nLaLZ8afm5V+ZKN1ag0N7LY/iTzO0kirzYH0TmXtPbCsDtwIgXr7++4RJrEDp4CvF8gF7uCXoTYW
Ux+2IRjHs68fsuRmV63HD0sxDjUdkZndTbjXo3oLvxc1wRqTJaP2B3cG88nKq3aMttrZ+W68fKov
CbrDQ1qrC2d98ScFxAyHT9EuRPGske0ylRZaHAfq1vgIWb84XNxspLyxsU8ZJJHRqWsTZJVw3dut
7PvUnJaeW34ARa1uFPHygTyqr8XMZ+UvsEEYPM6FIEXY+MY6q9KU06p6H//TkV88Yh6yu886ALKR
nckAq7i5bkJ6w42ad1TeUQrYEtt6F6AYHl6VPRjujn9KC4gz2XwIQzcEwqJk8LZEE2Dq3ZRAYGtf
Kaa3eEM72A8eluVN+/4sbeAwgfCjBZfm/3A+0SVeTYRukOPg+QKKh6muLCmB+MwOz1LiGcB5s/WG
09eYpTJiltXsffeEVORgh9FSn2naHXfawc+RNO7coLJmx/utQGv2vGZW9oq+q09erJKUZsD6eRcs
wwz+IaXaGftCKs8TDHrRPyKvSBFc1WNG/tw6qbnGBEbw+PWgF4gFOnISaaBeV5IMdvEH5hfVGZJp
j+2KE0vDXaAmk5ebAKRUqb83u9GFK08x3IXO7PdxFsR4a5nxi95HB7+HzocHQY7dPitDoC0LHoYZ
qiDnRaUWBomS57+MPvdTFkwUl91XJkl8RLs7Uvic5OXTbw8oUC7aC5c0D5duYtNKiVaVaXOW+6a1
HBPVvXzPMEyEpddwoVNhimQWnJdYL9g/6uJjqM60llImCyYxbjLO3VjZaLiVRaGMDWFSCJlOsDiU
uqat4pfFoWf4hPFLjqlDv7G/MAi6JLKAOt6OChTyAdIIpiIEzy6iGD3A8xShP5vYQCRbuG5BPPEx
2UIKDt8Dl/AS6OupN74IH8R3qLYAkgVVeCvrbOYv6VBlKrY76k5QrjSLkscwfOgdQNb7wMZ7KXm+
uswPiCFNC2vqfZrc5CBWWpdmxN9NH+UgVKOWOqBJayVptS5UUiwD3Zba6VTzE9YurXj+9eNBomXQ
4S/bULwpDSfTZ++Pad7iVMPZG95h4yKH8dCvmU5RO7smHTTrGUtJSwlGxyICmafQ3xv5XDVr8ash
uapY/tQdBw52jRlOVmChVa2RYqa3VwpqHBaZ9oKw6ZDVDmI3OHYMmq43kpeYJeSb4LCUA6Hh+9Mt
bzMzqIUS64hGWQorRrGHCcDAeZLAMmZslExcaNjz8nJF6Ixok7pqYNx9c+mkZswPznHTOfgRFLPM
BlQVEj7E8sRuNvHjJxmoy0OKJUgN/zbzA8GbGZYtYMVIUmxHMLt2c3FZgGvpjd6FJvhz7c9FvxCX
uoYvigArpH2b+7mzBvYJ/8XNa6lgKjnnFiCzFpsGhJMROoUqlHzoGs2HuQFGFTprenSbqB4vFFcU
0pwMGerTM7Qm59Gt5zr5cGjXNtHTfRrmLRmerSH+QfaXk/Qgw81u9FqGq+WuCmjwBnQWbMeEUTsN
meEWUlzK4aUBpo6R4mYzyiNT4vGzLPjY/h67ky3MCKm8CmK4daVSbjdGBt/na+TgAxbVI73oTRF8
yAaEc1Ue/i3FpYt6m2hdO9+/6xIYdwgPKxFmJ1X++sxQase2vIWSU9v6E+wrEwdJ86AgyIFXITfs
Z86USlrNttS5gxmYWRzT6PRS/Ts+EqmkgWpktiiLYzTSb4if8MeVq4w8lE8WHi0xWzyf+rkbxiID
ab7Qu2os17tqvEsnDsgs4OzJVEpwFT7/cchuRQKJR7DHI6e5G5HGRyzyHgz/eRMvSOd3rqOORN2z
lFJplcadzg9e+ETJVgOcx1RSn6FwTUYRlzi4nzjdGrxf+r8h/T1B09YKm4fDxOmhtIriepcY+fFU
NN+iSln2RUvyOi0pug9sADWb9RFAVMPzPBdNCapibnvxp4qZOOT95KAeZ2AQRNfwaj/lgvnkVqt7
olidyPIG2UHa+5TJkkaElIJ21+Zr/CBxIfm2wE1RubQ7OqUYruOUKpIYO86NPmo/v/pN5LFEB7rD
UKr7g7JBLaXEhS9KAK4XKhFybw6RMW7t5JKhan7yYI4g8Eu4cTfWLIeWXyv6VO6PYZRj6HS1Uoi1
ejWsfEGmnXMTqMUuzCcCsDvVEAq08HDtEQ9n3nzmUga56xMxRFPLz3l4orwEkq6UYuHxNEEwZ0/D
rlDtQqNLLPqsPLdNU8uLuV2beDf5gN8/rIFa0HUFjIFJYGm3gUEi7fddALZGN55SWr+R/cKRoIUh
+R3BPkBVu2Ti4dwnYVakyKEMN/c6Uxxvg5TflW2zdXmC1+9qa0I60rPEWPKIv8VH4v09xTkb8L3C
sKM3ZCGcbuuRD01apjUjkFo1V7nA+5aYNOpbZyE7xdvC68Ni9JJqvtUmYfHW/5swMXBupCsn1rsD
l7bOkyZxZrvCzU1yCCNY/mnSsR0Roz0GCrDD/EfRE4Anc0Mkv7ijw1zP027YA3J+Q4pT4Ww0X1qB
zZqasbI7KZcev2kA5BPadXCSeTMQcAfRk+B0LVraDU+bgdzJGxlZ2jE06EynGlfFU8Ex/x3s4HtM
UC2fhkxN1vlOGxJJd71SFUK1yq24VdW21FcT+K2aW72c3QmU+A4lQr9iXZ7LSwjxaYYT9CuSLPyW
F9d8mfC5PlXH1meB3yk9barJbSXa1wdJG21BMJ8fMvmAGrOc1ftTLlO47TQhVYVFlxyLn12HvYIs
sgNMtXPtdNNBtX1j9gJRtt+1cvupjU9meJEasm8U6TLpLhGMcrsYwapE0dz4XYOAqO0lXsrjBzSS
RvsOn63WzvX5HFdTqIwkh9lmRAUP4PztmfFFVMzFXTWEqnjsdAIIy/NAIRMnk5tMlT+PoM0CWzH5
33O0+RzfLQjkrALiX/kU4fD8jZsllCUGFaNIPbmWSARkHRHTzwRe+yD9T+m27B1mZInueXHxGWwV
qeg6EkiFAZg+OFSYOC1oE6gN7SJATh4PhkbOMI65TmogXXHlmwpIqPoJoPfOnNzsdR0m8MYLQM9A
gusCGBPXdf07YCymTE0/S2clTeQqk8WCYFSP47qsQXl1NGGNl4yEhGZXZ6W8XeF0FdjfNriac3UV
nbtYq1BWbyOFWyfT1Y3cjn2A5jhEXLu0f3MOGdyGEaqVnNhlbF61Oa3DbjUGFSiAOYGgM/vOB8UM
uPLqVUhsDorgoayQ7OJC88Cj1zbBSq+lnEIOJHlwUnBve89e2SvVE8UxQKRQEIuQM6y1PT50jQ/a
0sNZbHfzmz+UHRNZa5oyvQ7ykQALW9lN8KtkypIyJcHKbHtmILfo1A0Dgy8//SpNrpCGMi8hr87u
WH+o1z2SS8wR7x0Dr4mllVptnC/d900jvTJ2GBFSwp57RXLB6Zi0bq0DY1nSkzSoMmn4INIdGIQp
ZX6b+44XsfeTKVA6II1WqrnUPv/uTapU7b6RMkPS6c6IJxJacAVDPJoJdBP+YYvM++XGikvC7CY5
vnejNal6bxne8D3kU0iCrUUNZIYArYqsbgvMjWdsu43Fzkn15yAEVaFSEhgFc/JK75LCkVPDYLpE
vEhQ/iAP/MmwEKKhg7oBf0vxXrDVlRgzZBVKIWszKtqkAOYl3DSFS5wZ51aM/8QguR8iNSjD1HR3
WcNUaurbWcLj+E7zMNeHUijbsZf47Z4TYG2gZwXeftFq3Lh+4NASA1W/LQbpnsVdAPulxqzOIHaL
AU5OKI07U64a5WH7N8a9VHRudhp0fvLmnwuC4l9dImAfSfYJQegHpJaBnalhBaNjNUQfwq4LEnTF
JSQNaJFCH2Ej2mvNC9fUVMIjrXPpq4O37I+bOsfpfCN2bHu3DafNad5jMvXDdf0SyVpwyJ+5bUBv
umVQhB2M2Rx6LhItJ6Q4SN35Ao6jp0USQ1RhStywZri0Ul9MMt+SDWVRIw766zxQUwb/ivlDuDNM
pXqkGm8fDfz7kG2maMMaP45OaVPPtDYwQSJ718VVnegvlZGdkCPZXxmjumXPEYi6ChkRTpY+sCPq
gfm2c7bxh4OTZFX7n+pEJK1TtSDWVpE0znB+oOcFEafhr0t4Y5hGfcbcvTPpavSOxRoWRDoJ0zGs
8FXay0aQZjhGCo0+2aY4wA8lDtjdHQYsWx05ZvpDBcz5/5wK1/NkL9xcNMfIdh0FOt6v/5hl0+Wh
XyYcPSCDthNL8HRtNZQlICyAPj9qRGbBZ1JWFfmG2Cj/kz9fpZYDu5CFCq8FINJkMOPANLTy1yvJ
x1+e+PTQ7TtJXR+3xxqG0put76K6/pYfZOFXTeLQ4C6CGHe72dxcjvzdn9CxhLDIasR1AuM8LR/n
LEhnEpGDbeLF3QfMbYrOqbvoVweXmUYU0E4f6LQUkuXbpKGhgIgtFRZLWGYsiN9GfFluhHT4LNxh
ko61pzKcGBS1Rpw5MLnviYJExjY+ihGsLRkbWrNPeQ+kBjJ0+NODdZ+2qFNjIts3G4aDWiYROkRQ
lV7nbzCfW5VvkqnVwQe/yZZd2dQQuWjwVDu8ePlKlBr5xGq4Kn5tp3YrdLjx35oyuMTE6cTtfv7/
Kf8lgG2jP4S62nSf7nvxp4LVyA2v0hmhlUUCHZaOgxQ//SBW96jsqcwzZmfhexjt6P4CsW0v6MYg
PSHBfXlI6JebbYKM2BUDO1Pq4MaCiDf62vnX12Ez+WkPX23nPwXSy3n3Arx4kU+qXnw1wfHs4wED
EzG5cP9sHEGU6I/5nq/2FLkLub5vzFVptBu5vp+5inoBCA/2x4d1tm3yDs+GIPgk7GcQSfXRCiF7
7pr0IAr2sYUw9+biyobH+r77SORK+/ABWN5KPXSv9FhbM/X0u+4M3YVVSMB/dOchm8Aazl3i3DOh
eD3D2HlWEsHPScSl7jy2HNSL0tlM9nZtXU2znBZYdYIMsCl3vtlcDX2m4xqlnboOWgJPrFsRFDTN
ekS/d8VYzWzYa+AJj+wMs75uoVNYCWgM6No8ohk3RezfW7+XsxO/iYAvhWEM+7XKdcQf5ICNGdPP
EXnOejJr7GIjhce1mGJE8xp+sFl7qSUqnRzGq1Q7joiFLcQReN3sd5X+kNcdV8f0CGiLiRz7jjjm
/UmvCRIP+8JtK4mQo6rN0d3F9GYDyUMMqR9WxzPVoLUWXtJFdeMRZKpxxbdwWt2WREpLYajZU63z
eyAw7V8GMrtgvqxr9514mwzUhhz5rG6yqhTe4DVI+Al7psm/elFMVDTmpMru6qlwvBRIcNHecteI
5uWMYLB46xkDUChMapvW1i9+ONGmZAmmaLVUlRtk/sxp38SG4QuB9v3A7K7605iKU5qhRGbRl2BN
XIvQ7PVzWdyKdFvjOziqDE83OnQb8sNytgVzO1Ifl2RfCjzFINLT0Bv1Q0FaVTZCheOytaa4eag/
y9+pk+9Oy04iMBnn9E7HLFpn6IG0QQ8EgHakaeKt4kaSfBV47Cfrc/npgoULUrDpl4VC8EMhQfFO
+x0I6YJJafsKliYG7qbG5IjSCExkq1vGPgKu9cfgyCNeXs9rR4boEtuoviidW0rZVMz3fBXHsxSV
Z8OeNa4K+izppfTnZxCLvpb0/7vnA3iVo+pUfpW6jFNkOJn1oZo14xJpVdOGLL0KH5xtuwviBo6h
mxfEcehyuKUyEt0NIF+IxYR5HSpd/vHctqnFsVo7gL0dRgIICL4fKvhgGFoZB55UDjarcE+tWft/
CX2SYGrR/fHybzMVDJdaMtckG7sxn5qX5iW2o+oxLBNFEghFsmJ57JXSnnQqGF5C5KegEuMmEZ4L
cyw2KFl3Qe2kpVAfdj6qup7KUjiZ6QGXDvBE+7wfh4pamtCbLhFic18SVIXh612P4s0bFAOZNVj0
AiHd3mqpdKRGk524+YLqkPJ/EaKqIT5QNs+W3Q4wQRJoGSwCyBYuc09hlgJZnTYjKz04EXCDGdvt
KUlMmer6RtXUgZ04oYlXnGA5+960uqm95qzpE+JbBiXkoRP3g42qBq8Ck6CeGh6drY7BEcI/Y1+M
yLNBO/YyZywhWAHq+omw0K6Dksyvql3xHj1sum7mzgzsOJKCaYWmdLkpyOMvdYiev/LyRxTTmT//
SsHn4b6qVAptdNcj2a1JCzIr8V9fSTvQ04Kfm5SHYiUMNWOh53CiYq8zxdsD9TP6+ntnw0gNhrhU
dP7FHNa+GJOynZoU8KDWzP0ZfRkBhCoDshTOcz0zmIy23NX/vlHtEVHJlBRK1mjvl2KnsQ9NzGPY
p+c9gwctAIrwi4ooAZur0/tMlUhi27Ip9VJP0R40GjGVWw1rHgx5NYC2kn2I3eC018b3XfFWo0lW
yMACZK+O63nriPa/MK2m3spi/sxCPYdVhY6+BZZ/mYstjCfg9ex1uit1UhxGHA20HHGMqWWDmyBS
2+8C7/FRwdYJg351M7qR+uLshWnbT5MjN0YZ6mHcYSwZ+zLt5RA9vQReA0+m7puQ8RB1CbOXgjVj
ISUY2o9WJImvwWbXigwV/ka2i1+IANpH5245Xm69bXh1NmJyKvDtXK777EL6WJDqlVTf8xo9BHeo
tG8F0TkNHmt+MM6IZQE/lV7PQ0lf4r0KKt0HHOXx2VubESWlkATPTTwaw+qX0tW/TA2bMrqOpzDV
O9jRdmGr6yPnPN/MGiK+Ax8B1yh71olZlw9Sb0ruRz/Zh3TT05nTp4lfq/ctHgfo3Z60staFIGCN
xZukK2pEF5kbvV9kMSmKKW1JLLnGun/G5LaRwxUlN1W5MRRX9odNiaOzH/G8nlGC6JgXRfeRHl0F
gsuS/X6ke4ec3xa7EGqOOwQpHJDu2LmH5pQh+fISukLWeVVz0hX7dDEUvHEdh5p1ZDheaIupi4CF
D4R/iHwNQV491WIlAI/P+Kyuy28xRO6rCvkC7cRFpDHhyaLdVXeASZ2dpzlYBlgfubi9ErE3zN5y
waNcebifIQYgEjs/71kV5CazfEIhAyCKrX7fh7Fe66qtMy4eaJDqA7gSnFO3drQ2TfZqLBDktWs4
YbQmeBW2j4mNIhsQcsMULZJ8w2HpjBIqigqzkeYA55JNYWJpgCya9WdLdYsXrv3ttefC5uTRAmXw
ysNGzY7JqG76m1HbX7u4SrLGvd3k2NOF/eEfggmH8igQoL8No/BuI1kk37xs1V2LHrS30C+zO3hT
x7cyvGFoVttjUp/GJ2fOy39mK4OBPtkE93N7K83uBF2BI2XAcq8JucvY4Jfl8xts69Vie/DVH+EM
+V4e/OPGZEq1HRKNAw5Yhtz6waxC8sQ2jW5x9pMGdHL3OZcsR/dz9Vr4U9RSMSXBcE6zyxNP7uC4
mcF7xTtMrd1s1fB4/Yc1Ir05GONlJ3xhA76oQwFoBI0YscOPQr7RhzvWd7vd7310XYT/ZehNTQkt
IP7E96oKPamWSxeqPJlQfxOzW3Qh1ShlLpVLccJcB3BEuZSBZHVp096OZYxUEJVAiR6B4TKLiRb5
OvWn9+wowwVmNyrBdUQ9vD8fUvTeEVwEwL/9s5YggqI7XWd/z3gDXERzL3EoNbAzR4fD7d1qWdPy
w47CNrtU6AP54Ptut9JkuR+mtW0jHqeUA/XaRMUJ5RgdoaPEEktvOty7wHx5WWUtIT8tBqhG9Qfc
LvJgbezUUlGFcz/3+JKurDQ/H9nhYWDyWvGuC12jcDVyFLr/K5fFRYpd6hX7e16J5jo0LjQvSiiA
lq7sYf8zrDyDwqPsYqn7EcOjvIyO0+co3DLP/u/tC+ohFjcZqh6/aV7q2d0Bh7cDsVC4Y9DetUd3
i+Vu6EzBmgOanBhTRZiKtL1H7EFDXQA5isDcnu7XYTzAzHZ9jfjC+g4Dt9KtPfiWNkcYyOyBofrq
/mZnN80nJ9fmkPUtVot/E2chx9j9fGeeP3E1h9PB4g6ofdrKi8IynTF4ed1AR+3sS34sIwWNIK2F
SI8qIsUDvguWjDu3bk2GsNEJS2UHox3lNiBeE4N+WU9rsLbnabHFwGqlDW4tf8EvuECQ2K1V6q/q
vRQxxu/Y2q9zyxlFGQzqxsOcGGZQ/4egmOCle6jimD80Mxk3ZVa/0aOVU8eRXi5rTDJl0J+qmW27
Kimhi2NAiFyrqqh1gY8/QxpPsTE7lviaH7ekgcmrFWevtXC/DV7UaliGmM3992mtmra7udO22WtF
rFlxbDWo/tMaMH4yZevDnP/BZO4/hXrrIJK1GYQ/FhcZ+5QgYTcq1rqTmW8HbTK42f9myqp3l7ys
leDe8X3e8V421ohY71HoDN/dJ/5rdvwfe567wFsCL4CaJUYg9YW5uklR3G5SkP2HfiiIn7hEm1Mx
lEz2rqPHYUdZv5sDWU13gAXZyNqM8rtsSUlrfTzRZXPtWBPfacrtmJMeMkiXkIzFYtf/H3CE4l3P
RPZdVWSDrmzzcDwcdxUNcpDp0FX8YXXwjvt2VI1JDWzT2Dz9S+Zq195qJ9/C4Z95We6ppuFvHUX5
Jl7D6A8Sh6/8tsqcZxQrHN9Ap9dpwyxWUsfBBkCKCnpZT11xTnEgPEfAXUmBKAxdd3jzXfoEySP7
vFZxkf9ZLShCVCxv44P4+FBABNEthy+t07h6I71S24WTGg7AZaxDVncB2fUBV2ywv0m692oHDBI9
slWrnK0za5A+gFkLozQvS0WarekodZfvN1+69hj/15Abb2+ZksZh6YxCDatsEohoU44qhMIUh5SA
It5mTCaCwNwHAeztdhs1G4hjgZeZzO+WEbqnSf2X1u1s9hRRqkqJVnaMD9gJ6pPo5i8pwTk2SBY5
130AIZlirxCsI2t1nQXcFHzI4EJGj89aHm5PB/npyIcubWWy7dgwupfDGLiXmc67dPl5v8vdnkBa
z+2UZWteZIeSK9M4bbg49jzWGfVmlUPZ/pKvnyHhGNIsr3uuvrgSuEhf7xADsNiL37LsaYSpRG7C
L34mudJiQAjaoXmPRQJiL5NNkyxpLELxmJGl68etXjxIiPFDDECXkS2beXiAOjvRkb1Ik6v45ANf
X1Tjp7dWWKqVd8ZP4nSLBCkJH8yXTwGzd2CVrPVhlheCdheF8959RwlGmj8OAdm/mi6SddycEpeg
87QseS3H/97gky75a7OWHUBKQ9B5LpFGtEWmAQH8VngOjqoR2W3sACuARnzGspJy1Mb1CvuNbSmr
4bx5vXt+XrOZoqxAjjdiIHcPAcQCUZ4lHw9dTqssUKa08/rwHMIImd+VyyxL632NTdf6fw95NUip
UcAokY8TMs2pImshgo1VRrFk0i7MA9tBQObusIV7twlq7iC70lh8Bz0bHi/Ov6Zq4Dc+JKRkpZlU
RMZ74GxSkoq9WRyZkJVkhDYFoZ11hJeKq54OftuUf7l/Czef756mKaManyOtiInrC5bgdpr4Bzu8
4bD7YnmtDKOhOp2YxJ/pV1gy8KkWo6ydnypqTrS6K7W/DPR7esx5vPPTAoiTiX68IRkP7W/IAJLW
95PY3Vv86+KetobeyrCiK36eSa7Ix59Nwb2CGZEF2A6fYuccdZm7GiXFjUYxCBrOvOQLCZKazm8D
+TgyIG/SveRipwIgDnOlGkLsdCm06FI+pMo4nIrGYq4EoFfnbjDxUetH/UqzTUaFAyHsfXEHUgq/
I88tBumCwDp32tJbUXz+bY/rtoqS0hDpspNSMGjSoxdI66e+sKjTIMoWviyX0c5o4VYbCGsDexdO
lUmaWhjjIQsKC1Hp49t1h176Oa+i0dXGjnii7iRNjFl+hnzvYGYKdbhWI7HFMF6rbByqJ0p95w7E
L4n4/dMhKzVVz68YHJOVT5jL5/IsxsWU4Ljw6vUGQVZu5GjliY3KYiXBIh0Rspfdu0rrQDuHkJNB
OtEB8/TEq4dNVvAxaoOElixIHUOJr5EOZUlJV+Cyt3037RcrtQQ5tUIru6SJNAKIRSKXx6pKuDZT
+dA8T49WDBo+qJCB7A2ZJMbxccbidBcyJxP4XgEsxzw8bvWpp1Qds+XLiOSf7JtFTwK1WSfvjtg+
wSz2xCXM+yfYuRNWKMj8uXaNNYp7d8+2JrT3suYrCbrYM9ixBX3FxgpWZhwsaDLwrtb/65kkIpd5
2TCdbU4mDPM0D/EUHUc7teoXi+xh+ore224R7uCT/5VbBHtyQwmaTc4w8jpcqO5TUbRk6XEwtuVT
FxZfDWqCDmDAR/7fcxinMDv6Z4ZA9mgVWAOyzWR25+kNmfvfxmyBDPNbAMn/9szmDT00nvbZQZHN
vOpmfIJQMOmEC0gnIHd6sXZym0IhNfQLSqFX/57M2KlA9mGW86/MuSPjwIQfcZZW4ImimxjiW3+k
zecWRlUXBhyQOr1RxBau0d3mN+TosYAi1AzNwLHgXjGtpn8Rh+/0aZFkSUYfxoU6N2dyDZRajdmN
/0alKFVP4Pnyt3Voe1B8Uuiz6wexnskKHe8GtfMe7eEF3Wo/fm7hmfe3IMo7JnbuUDNRf8Om5TCH
SEtOzn4sKncixEnfVbCk0UCCOJPWhmbNsg3u3GneKRllKyFPC+UGLRYoJLoTVSc56/xgMkIuTX1A
6zlwvlWoPrYlK58cRorgywH1gMMd77w2vnyL6yjdVUEI5Ti+Pl4SZW3lOX4XV3inTew42QHkABin
qmvOP4gBMA9FzvuusNWCw6X2CKx4EJNT1+YIxrYtLKRTVZbW7TROgCMdwWJuLg6dQORRyYGI9gYp
S8bqGlILjDp+toqIs5BLGJb6H/8/W4LPFaAKvHs7pvr05OCluD4LOhJetOZo9xap5rmmbkvW3Hgp
MAA7gOjd8k678YJOrRprURUHZSfdPRyPGO9sh3Kbi++pQo53hPciQ0SUTrKp5FVa14cH3d8mS7SS
R0IGB3occxcH7DuZBlG0OFF7jNYGkinpmq0Sy5UOGS6AlaEqCwBWsEkP1/zNAoIpAmKJ+QuV6IGy
hkYnST5MGAoModmoEGfDmIj87raYL19uECt7Wdya02XLvOH2ofqj/JQWmqpi0PIdqXnOt6OIohe+
dg3IY9fuFEXAkrsWecBDpD666Tr4iZSb0tmY7ozkrdXL04BPXoChd+ARdj5C8VwYKLzf90w9r8O4
zssjX3E8X5mm2zsKCDos1pXuIzPIDSLR8Pr4e2boIV0s8vgzuOK9/bKH+7DQNTfse6NRfhzDYUOC
2RMutVLYdug+5pxCRoIGLs2XUCc8Y0RH9d5GinthETmjICSlD90S5bjop5I8p/N9d25XpYVV5p9I
hH8/ETW1knbmjrZdINVhGT7E4HbUEPf/BlCth3l962+hd4oelPOGtAIIYKI42voHufDSiQ7z6YMs
FBvtVEox0tNC/26BwjCeq2/oXFIhyj5wKYF4fcOGnr4WwtlKoJcpKg6+z2/mc2mQaG4Zj/JDQwaH
jPlHZd5XFXK5B/q9SXa1E+Mx+vmscR2rrE64kQDHcSKPGBYEAcGEW1XL8TqxbE1uHrOxKrtqPLdr
lhO6ffMPHsO2HQWfqK9uLK4FdMmMfVP1THOb6x8lCrxCThqajYnmvIQpXUgnXM/Gw5DBs7dzkvan
SpGBKC5Xq/5A8elGSYtmDsfAwGa31+51Df4b8iG1rkTKiMDeEU8v5DoGlyj7eejY7lxQrS83JbDf
ZTeaVSPwD2PaRMzcN5jXW9aXDVo3FKLbqLlJJ5kN0rxfoKzGG5bH80FSsGcgdRiptOSgMFRMU5Ti
QhLqrI3WFj/lAcKDkkgnZhrqNwThVQ1BPqCn/dRyTyG0yLIfU5PGd4PFbwMmttlWDo66mLIUFZ81
vl5VG+lqvsNv02MaFi+D9TRkRRh3clegPkB2/q/+/J+ZTKsRIwB3zA556yJhsU5huT5v17kF0dmI
K9RAYGXF0vbw16qIoDr3j1sqK/7oakevkDgLnNlb5nTeZUwH/cmKb06H3mxx81s4g2xGiKM9kpx5
N29Jko9exSSlmeQFBPH81M9ORGkzCmrskR34HII2uSZR5QN50N4J8RPWpp6c8psD0t8nZsSSJ1P+
uMxz27cMQMncpoV+SX56fYeApaSkMNj+pLUNgYwM2DKxgxGfn8s48SD0dhxxXScc2uIDJLGiD+To
0xSFrNZmsyI/FzUR5QaNbsuZXEAKTHlBGBhtqY3gxJA5kB5MOfIw2XSM2uzdZ9D6ySwKXquFJ2CQ
zVQ7pTXVbPSBDKcJL24BulxeqbO8amGIXukUZOP5YAcdFiYyOEmI/w8PgNgO/nHW/MgXgvggL1C7
vmA6o2eJPT5y2g0BlPnI+TzRf8YDiv6PnP/IbUlGxBjfnDENZLhmR29sWC2i16Tfp6fsDKDg0iAY
gr25cxiw9wNdc4x5cPFTBprcQFmzXO4DIuZZov1jjhqc1n1mkXZvzgGFbMva4deexyNiInhtMaCj
oh47NglzDHTkJZYcIpcb1FxdcZC+yJluqkAMRVIuVYGizia8hBtGPlrL6Jy0Y72aSfumbhg9tBwP
p4grgwky070H0J3eEvi99mywzzLQGk6ZqXgni84kypmXRDj/kVmNoQJQhL/L/VIxsQ4tV+dfWoS5
i7wTJGAb/XW46lsvI6K7glTEbwnZKi47G3jBksyLePhc8q94roxgF1WuznoG6HLl8KEOmlUhKQBL
Holul7p+OCxi3KZgkVKygCzKnwtBmEOQi0gjOpnBcTUIQ2DCtRawKJ3w8N/aa6Um+IJL2qfehipg
+5XdN3feJ06MvnIkk9udeEn+0ZSuDhlcjQK01n3kdK3ZppLpRWD093m/zlu/lqhljzpTgngstGjz
7Or7+AkjH+9BdiOz0ffAjmu1QZ3W7MRTYDeKbIqCunw57iiJBwtAgaFLLa7w7TkHZceSXPsJ6XWG
qZ8/7PB+bHtkPcK/ES0DbvR27SLo+UY+LCTEoyRAaHDNuedRlKoGZyAqBmyyiDk7AunDKLGjlro1
b3QESNJ9URIz8ZClUk94QGjV3un8QJ/5eW74e/nB3Ku0qhGnyb83jgBPFrOoI5NhhiCe2bqgt5aY
gQfdM4g+dfWZKksUtbWzPqC1CHI/gLklY+VRTlEFpxU+0P3fFmpia5swZzwE7ISonTOsJeKgqWaB
PE9uoVIBihRUyVusd0SFw1vlwFsw4f0pu5s5c0Dd5qlRHHZ71P+vi90Bsqehx7Hw8y3+QIFO3MUZ
zYjSL+2FLxSDHiTfavk9/VCxriYR8lnLRN9UDZVViDhnNJi6Q6XwTSD21zDKLjYinel9vk0Txaa8
ovgR9yQ5MEOqgC3KW9j7MIp2/wOb+U0TKFHNbp8eL4jbf81lwYwhMQLiFRdNQ4Nshx7+VE28fH+f
Gy0LD1O6bxUSN+Jkzl46qIfNBRgMg+klZhdnVlwYMLOISC58kqZYTXYBjX/MThXBqmeJMjxl2OQk
D2IDr+HJVyQRSXE1iHRcaqF0JPpl2QdJaA5kHIVawfUktrxhlvUErVVi1Mkmzi51fgE2RvzZLZje
fwcnLlawYLqqpWO8jGqU6GEDqxV/ZwiVJSpZklXMPV9GbDdv8ADxaQ9No55LlQntTa6CINjkXjDr
SN6H5L3wipNt/kV/TjY1GycBeQt5xEt3tdzK6sWfz2JTGdHhcRZWjA4zRwUzNiElP10bKmJBVVBn
Fx0Xi2JUPV016kKVyeun4v0PoX+o6mymqSOqIlTLeptbake1fWw9VrY8DGNPhNTDHkn8ryBNKxph
rrx73DvzYjirSo7VPCLcCewNQMPM5ttmIdSy7DxtpJx+uaiE/NCv0Me/v0l3Gwt2v+Nqw1i+t0a6
J7mrMoMiZhTSdf5EW3eMfw6QwtteHAorHXPGdBXUrThZWwFZirpmleiblOcVz1+MAw+hCKDoD98o
folaxYOdW9rddueUa488o+z+shRLDhYkJdpA+Jl4IVtd84M20cZ+nUpKScKB7CgSlP290J41unBe
S0OzhYJiUGz7eZnDW9/nMe1neZf8faM+ATkj4SFIMi3LH/vl9FXWIoIxyoh2Kl4H0eus6BWnUb7T
UHblR8XtIvs5OSsZ0F4MdqxkoQ5H+c316dVFc8XzllTt14fqLGSYBD2FF4AhH+/mMJvTI7HdLGEE
Kc+IJsUPwqS5F7PG9fjCX/e3RFPvj/jAjuncTYP7lZ2vpWrZmjgm9m3NLlrFq/GDLyW1WT7I8iIS
qCz3JFW72UApE3wouXUKoIIjEDduU7Eu5mC6pYfO/xuEtR2K0f52FXE6vvmKibfDy9n6tOy1pJGe
Ej6Geahq/XOAdcC0NnlNMAZBhT87pMqgIAowzCgvTx23Ew+ekAC0xBxL5LGPV3D47B2h+undIyq9
hmwmFjmxAvc4xoWESqthLUEYsoSGsJVytOwiPUYputQgjOeH09lgU4yDyu7cKzXY4USj1y2z3pnH
uBO/u4g/VQ0lPRQ9viuNIGjCSNpHOZbdNs67oX3ntBOOLOfHTCo3gIJ93klCjijUrKMtZVqwmCX5
8gG5ZpOmiyYn0XNZSZwwNZOMX4+ZLAItBqpwX3E1ntur6JAzo+yKYvUqfATN5FNKz8VP+N1HDBu1
ju40FbG6F5BPLNyMgYTkWpXQhMQWDYfb53pf+uwvAO2zZrRa0DgNF1S/FT6DGCXF9HscLIzr8ZGV
2RuPzjACIXhmSWd7kwY04M7zhchMMiuCZ7c3tBZNSRl11+OA1riUP8i6AqmirhNyJntTHSOkOaLY
kgKZaLwGvf0A6LfpTCIekXUfjTTjan7MTl9KkHRFi6MU2UVJkI5Aov9yToe7TdZLqglsyw4X916s
Eq15ATPZmi2TsH8xvExpK/9VRrnuZeJYqB9IiihX6B1inh6qls1pNP8Bmw85TP3YBYAiwZTrAPNm
0aNpZisx23HnEg9A+ZuBDEu0lyrio3v2Xb9J/T0IYdHPC96dREjN2E/KUrzEBVIlHPp8AwXQIt1e
OEAuDNB2sNEZfmylAOonJc+f1R3c4Cxf7nfOFBue4ilXwv4rQyo1EgPn1K6+458XqLZEfya3aPcU
gWe1kjhG8m23U5v/t8HG0blMbUnkYH/EM3FCAlYIDb37UybJOt9T5ZSSvWjsrwMP0hx8RqgAMfeY
3XoEX7wytneznqju4EzcF8DJgr1qMR3IHoGK+ISzg/PLBZbLiyFBKk5cpv/KKSX39s1WaujnfsLs
NGOIimf/rhiblaHCF9h7CWl69POanO7qNIMAmVyi1OWBMHu4Vi5/sE3k/Hroyp4OH9SKI5cp+NZl
XxMORIql/Ms+pKEUjxekVugjS9p8MY1O4drC6LbBZlpFywD4NcH4SvY/CsjQwBBim69T3n4TbR9y
iTdJHQ69NWPoBtuDn3ZwDsjBihwbQAyXmUE+tTbCy+hiSfhuahoJi3HIT7iulKu1YjHwnTzLtuIr
Jl2DKTrI0OvXnIlpvFNq7+JKyASPyKfQNd+Kek4UwmXj+64XloOixqlOJvQzzJj3UJQ7iYZxnReD
6kwMTo3moINfkuMwqRR5ruGgxNBchsAj+dUIwmOL+dZjsC7g9dBUu7lU7+dhfA0QaKxEiu3oejIq
JktGtXHWpS/aF4ZN9dDKhrc8Q7R7SZx2ppPrWTuT29ZJRTT8RWeFmXoVonAh4uuKEYouoVj4izSt
QnQsohMBP+khxjbYpvIJmBuyT3E2ZaY5A3ae/IeF+X0hUiyFxscF1CyLV1TBM2bXl8QUw50cG4WD
c1RxSuzACyOsKbPBnWhKhN9TVGk9E7WVCsN4hKYi35hH5AZut0HFnvnMWoHdSG1n9wHBAxKD7YYm
DRfYg/DylP+hozdmbbblGKvZGF4QZsP4gre94epu1kCciSm+YKEm5xiyGa+Qf5WOtZ0h6oo5q1H+
TjXt+bdqgEukr6FTUdqpCNlctYuem64ERYDoIfb1vUfe+3dcZp3Q6kxAAru3vxYQYbXYlBkVdsZ4
+DJyOAhj9IHFlBZiXDK1VNQouDnvhk6XYIIJih5rksHgnyGv2MEn3jJRmWEcoLQlaU4umqUACOAQ
j6q99I9WVonYNXnE4YDEYwt3lEdhht7oXafXizul+t6DgB6G9j8S1+ZFFz0YferfhyWD7EWRo4GK
sxKAUrDzsoMES2tam/RmzshnxDwDKhK+ldo8yWqWfkdWt7SIN3BUBpWK04j4QFYqInc2glOsk+/0
jYdCAuVeHTXkc5f3qG6vw13girVY7ogDX1oRNxgojBDVLqiU0UV14THrsWLU/youw1UWLvnEesAH
Hznmje9DollZG924fsN0nTKbhqPo1nxHJJK6Gwru2mjNmPU4emubdqmpaqZTH4D8Aso3IkiYU7Vg
cNx2IvNktCxmniwiglNahMJpjoD8CWZ4kdS3qWGjLlEXNxm/PEpR81bON63bKaz+XCKRkCyoyCtl
tNWd8Lv9SpFV6IwldidE0r3Z+QceZMB5jhN2oBtDfS+P2moc3XNEN1soS1dLDveZ+rfNxuKkkyjo
pbBRfLpX7LF8ofpyWVz08+hxhHIfPOR+i68l580tyEgeBx+1WaQwXd36Xg3QwN5Q8zAGmNdC5R3R
cUJOC5qUQN6o50gXuC3HpFQY48q9RnWwqsvd8Y8pWlMlRoqtBD8V+5lne64nu7rIYf3ESOu/Rf/M
96XAAD8K0eoHE5shzQwokolRS2RjCuvxyLGW4gI6PKmNXrqecvqFZQms1mvmiwX98ti6CZBOe2r+
D/fvlIrVIyIqDhNAQ5z7XfO9prWlPWwrMPJqXR6P6MsTJUVIiibIxSWa1NUrZZAiEAIbfrocf0Sl
Ai5Mp3MUVgN9GU2ybyEiBrqHg5BNVHj6SDfXesmcNFHwypekMQlOAKjhWkRkYHyQ7jTckCRHvmwj
Bq561YAy5gRxcPUNlXtCTWBcZwvkJH8VfLluQsP7G8CHrWPb7rWgjJVrPZYL6kKt8soRpzzY/mjN
Zn1wN2PK52ziOlL3TrlRV9zjYzCGExBpTkL7Z479wzuz7Bm9Dg6PDI2YN/xxhd/Ln0jdlkO+0XLG
YkBUNsvuBrKBBKAZH0nB2SplbfIeFtazkz+yI1lu1yXkUZBHApDAI6xhBTaW1eOlanjR7N1PjHgA
dvsrPqtXANLi7SfOZTW5DmxYncK3HDKsWbTMsCf+YDY+ZXvZdAk9K1+oDfEXthZF4RlMja4ubs7b
yDMExn0qw7Q3kdulSrugx+jO89xuI2wMCMl5JPb82fo5VPbGOMzaZkAv8zwP9+TMW+iTcLmSkPij
5IW4xRD1aFmfymFK+Pe3jmWM6uI/wNxiF4fb58XlG2Om7tEZa/Hcsn9mrsIcV/jevn6rqtIoLUCA
FIFkwH0DFl1rgPhCbVUdUxgAMdfoGMRTQzU575CQPwXLk+O0wGrYjH3wtSdC1J0NiM+9vMZuM1uS
nU06kYk4yOEfSq8CF76NEmcrzkZ/fd8JP3s4qgEADBZqSfdK6vO3e3C5Vdfs9tq+DpdZSn32POfx
hWktHFsRUH9k5v/fm252WQVy1DpG4zm9LmutHaHzgq4MhxnC7XV+ArR2c2SnYLQQKmNPPNX9mNUF
pilexehCn/wZX0QZEegzPttup4dtCqisRSbD//1wEHCNdAM3QPCe78/8+lBEhD2raArxs7nSqpSB
AnE1qUiHc38aytWEMIFM1prJborFgZMiFkwCGUxSKXHSBEFCZfQEQloJyCUhanwzhVpQLE1wNooR
hRvZOFRH79lZVr1ax78FHINpColOBrvac/Am83FrYuiA+72a3hsVMazeHklSsjf7adzHpk3BnNeT
DOllmfLcBe+/synO5Gfw9KJpT0ZX2F1qb0UcFwkrXGdqHquaLKu1vYD2o0Z8VPe+ZdPPB5ujAHgu
iEDgTdTDfnqu2LOFAIu9j5XA+KOfj/kuNQtrzN+dPvakzT82Q3uaCzCFfGzKtavbZ66hrx9U4mgJ
SL8V9hJ634ss7ZTF4WrhuxP33keTgSTVpYMeE0Iy/rjgltXN74ECC7AwGDEUgCsLOm8ItIIrgdha
vGJbadO1bu8CWRuMTTsRJuZ9Y+QqsK+pjWtV0P8QagjNwBxvgynQvZLzhDs1TKVZd1TSUIDslCY4
OySgqnmo+7L6rqNRCx5yEyMn07SXz4pH7DnYTaMVLqXguk78kDfgKJZ6qpRx6hvRUw3Gwrem0Or1
nhGnury13rtJlCBylAQL7o0tg6RCpF2s8n5hbvMYWGcTyiJFfER2Y2/fqd6Vm3Dylf7RBrG1b/OP
wQvvx/i6LLHOOl46mjiWm9IULTcyoTtY3igz6dg/JCiKRNfdPXERpzQxU719e8cSAs6SbPXUQGkd
N1H8xQA5QxKf7QvejyTf5H/79MrYi6MfETS4/GkfDbnvVPtzTFizWQvb7qhtjz1t/N1qm/Ax92yq
mvmbSf/ri17T4gbU99qusnXmxlM02Nn4TjRm0JMHmJEV4mxVihSxl3yo5StKDe9gDrs8SnaQSHMg
Mx+tEKz40jJZ7hS/VKnWTM2LX7O4+xwqdj5RHKjEB1XEvCpJWjtKyfgk5EDx6ekUlwyaVcJXrU/o
GV5eIx/V21tl5JVceG9LLZ/RuKdlS0ZmsIuiWawRV9Pnu0PGQdFpuitr5+F+tWAuyEYpPZtHw1TM
n0uxs5qwpuHfFAjq72WaUEGOupYdHX32UH91J96qfUt9VdsIhhve0OVya+IcVjD+4cyfzxhgVIMt
UtLsqcDAbt0ujn1v7H0QjdPVq/I4xsfHbTapsMmho+ug85vDwFUtjWOSHPfSnZtZeReG+M/1SzwJ
jy+Wbre4vAk6jDDngxNImKAevRptDmTPmmeisQykNTHqBExyB3xzcjzg3wBaV8ZD5f6H52cceikb
1zD3t4YcmSOE2ITSOymA//k8crXHYwCbRUQYhnLt666NpG5hUtrPQJ1A9dSf48T1ldEmZJg1ihGz
UNAmdiybnbaGLnDzkjovzjNa5Ugl3YcTzutUOaVV/owil2iDJQotGADZIIs4Pxaf+n5GlINqbLYr
ETUBwOyuqhyBLk+9gjIEl7fFQAVWnfpU9fZ2O6IKhNOpClWeNYS0MboybIoSGocRZlGBZPDzc6hv
5kL3cvhwi7Vy5c7PlmV/ogrx/qcA8F8+vcth5WGiTfeoSiXS0EzBFHGvlxlnhfOdfD+4roQpvOsQ
b9rNdrP9iWwQmUtMt6qPTHQTZB3StNucM4HMAYC0TXbklcpkgoSjNN4n5rJRLS4VQEnIb63sLRTU
bI0nDdJmyHTYHHpp6vvlvK0X2n2gVbxvs3ruAxx0VQwy6N0yoOCrgnGNPdjqf1cJch1jQO+n6B/K
yt9tX28j4s1VuUJFXEayFnvmhFFqz76OPNP70eRreORns4yFRiPwrxzQKzpIqcZf7UMLHAWeapgF
+xY3qcCn3QAZs2P/tkPEnarZE2lD/iRMGDh6sY/DD5jRfLUvCcsMspry9Hlii84vxDabCsGMD5rE
ZnDRwnIDPUAuHcjE/kq8S4ebuUoOfdYrYCbeBFs7qzr1ffS7F8X42CWHLinYz0oQmaJ7e0lzZlRE
DPPxCKkRiXiv9omSaqr/XeZVB+hOGm60J4WUhO44MmCSrGk7SWbD3VFZfOc2hh+1SaFLJ/LWV8SS
BDAOFs+hJDF+dyvfieNeK2fi5RXKHjnuq9lIF2awn9JyOSGufSZoCjKzKazMNyL0jDavU8BgfbH0
ptkzbY9ABJDbuEX3KgXxzvHSCzSM6bRaKEvoSwPzz3mXzMKLe0SS7vusz88mC6jpT1noIW7VXKWA
94y72T1c5sGfh9t1CnxCznJ7q7cnr+C1nHIuEVOaBPmt3DiOCG/nr39zvodUixw/eeFG179yFmSu
ade2EWYzs5xgVVUaT9pX2K7gM3i3e7Y0PeSHNWbkYQa57fUxC1sv4kd2nlb5ooOZ84+DKmxYQjGD
7DFCricwHo61+gCxeThBo2PZkLI3YqaLR6dRFeKzDvHOLgK++RB0QwN0M8GEKksxwFg50VqG2T+i
wHJvTnduvmGPtXXVU8I6UIcz592w2ETiaJXTTD0jyKmMs3/PiAaU/obbpgMtDYwhs4Ru9tyiHcLR
RjIj0qUSsF7RBB3iKYI29OPcF5FFofOpK4BlYbtzzYe8UTQV0kGAzzYsBJee4IL5J4oradMyPgP0
1rtvF7+5VVdFf1SPLKtTo9W3dHPAxqLMqPbOWc9JX4ydDSelVJHoO0EkkeMS5IkkcPTeCpcXIGA2
aZHAgCM3WDZ64jxQ8H575xkqnguaXMZ2YuBfWgcEzIGuSUNPj7Oa/HJffeokU/kgY2//Bv7qeqnJ
d7xbhDPDr5rtoP3bLxUa7l5APPqOG3uo3fc3hupWeNeceSuDME3jnXBczE/T9ldd8zsjRSa2vVZi
t+kKGq6LIZsXJgTeWRiWHPHOHk4Wt+0F/AJUhp1m4AEtU0H8+4d4rC4vqsr6p8K8NfIinP+06JU0
OuSQX7MKZy0jFE6sfuC0WIKYQI6u2ENCSr6OG2IORjxWOZs9Ug9kb2kkjI7OIqVtLV3//UWsF6wM
GEkZFy7uy06ZWX1tz2qjjx2m0tdBQljFKgQ2G+mZpnCsUzNEuKuaysYDi7dV9i+UxxX70902fuxD
gT3RaTJp8EOr1jPTb31Hh3hKld5d/Ikb7G/E8Pi5OrcO48cBZISeZOjhaEeXh0P0gpEYaSHR0c9M
Az8btecA9o6Bc66oGJJsuZkP9ETj9hZM+nKEzZYcUK7UliTrsmtkeguRnL9ZTGgY21emJtiuk+Qh
AwItS81X44HAd3EVMuAFEUuKqNahOR6ShQHmLzTPLBTGNlctROHC0F7o3OzZ4x9nf/R3U+QlVw4/
kt6rGB1mXhN9hKweRKTTYDIvVwmjSo6Q2XFPpqkq34ZpwmTyBCGj8EEo9DPliLa6I9uX3lZsCqUe
OnHzj983cslP1szQgLw52MY2Rr3ntXsLPFB0D874z4g5cJwfg8CQ9vxsPkNfGLxeU5NTriTBE2Yd
t9HI+PA4047+Nu2dMshuhlTi6gK9oBu+57sNUDAdrksIAuq+mkwK1NUvTXNbhx+Wt61J2a7nMMqS
wW9MdZ/QtMasLIeUVqNElm8gygiDfiqqDFkWmOpE0Sj3GZdklUxtoU1EzbscxZsILQOx1lIpeSEo
+YwwqAoqx+GxgMwQColNpP28xCGEKTJvSNVynXvPrcmjJ6JGEDQBgNljug2jUl651K4XR22Xu4cj
O9DO0J3k9eU2ngK4A+Uj2hBer4sCvVqBt/ETaXi9K34VhbhBdbKiuD5IajBaz3tCXeIjwVaNcRWd
Rn4smkktq6jz4L6HiLwsijXq/FjIYrYoczTLNqQ6lqKIL95IkvtrLRGRRiuxIQLRfD/PUengCVpv
f7dfZ3/yxwSjcePIANm2TdhHZLVO3DIyBvd2/GCFs42ZdGvxqKaKvfw334EaMGPGMPQbatbed+Yw
e8e1+5imWxeFhDZrPEMCELS8EBRyJJ5dl3CI5S93lPCvtXmVMTSyHFfYypbL0Fqk5Uamo3tqVDf8
VxPrQHCIsgyO4uX3PxDEIYShIlAMsRk8PA4CqgKFsc9n4oKF5lsb9F1pO0cKvr/ZT8C+jF51ikzV
T3ksK5z3Af9vIzoJA9XtsoTwTiCOVNvwN9FLa4ivNvBrUZGJiDdiJtGz6zfwOVaOjtZNSe9sjcW+
PeQWnIxB7zOf4jAqVdRep2KcVXRK5eNHTo0B2wSquowwm9Sj4edu0nS5PoI6le6EemkiARHiaB87
gr1pgF0BhST7pCZlL8hb4FDua3kCnDyzICIpN5lI82DHtnsk9RhjyEsgVUs+g5wwCDBkdj/pFz/C
axotcmh8TAyjddrIf2q2i3hHw7n62iqIaDCk0BAQOH9qCOq534OV1/qLyRyc+euURk6/UJXM2pv4
rJghG3gPA1KC2OdtiddkKgnT+JAXuX4/cg5VuGQVRdJLk2KQdsJZiGHEwAFgSJoMhnRB5hzjzfFj
RYfLeNpxiqg+jKzuWBwL2ab2Qipwafaz2KxCDwHsRfyEoug6u/LFnD404ZSa/WdYMG5Ux6CSG+xe
lohxebiOSaXwMMqUY9z4VOs5IIekHlH+K/ebLW4dMjBccJTMonrKdGe02Ueq16MVoaAAtmWfTZ/b
BICEHanlZTcpiNuA55xLLRSSGEopbg/FLBuZ7/G5xgvUKFC9g/Dp+A27d5teilAb+ddqqLhwi2zJ
E6La9LN6M2flPwXSdNO2T4+NE0iUtilX12LnpH11Xm/DEucwDJhXII3MeD/5aBkfdUhUgXb+waAC
LPSHxHaciuK0TQKxpBrWuP6VZUjcSVV5LI+B2U1CFTOVd8qzc1V91udIDLr19+d5idkhFnJN2lSS
Zzo1N/qTfMQNExoDgwbXMCwe8WxAjpDaZOetMuoWDjcHmsCD7vbT5FoS5xuE8ecBbjF9duDLud2m
LtFmcd98SN0QqQrMyu8+h7ROVUFduximuGod8o3o8g9mzjPbuotpzg62APMO+9r65IEZ4VNDcH3S
LgfLo7cLgn2ynfk70P9CRSUB9nuMk/5Pw5fm8wqK6WcyYXPF5XlF0VODRa0P/z4/APmSBPEWN5kj
mq7uRVgfxV+SXgjx+XLBR8uCsNPOEUjrUeMeIUz3FEfnxQjk5/lWWCe7LzPyYe/DhWS6SZRGWX0G
ThzLH5LWHgbckYfZ9RYbdOWZQGHLbejZnKVafWZuFzYFu1PgfCuutsXKVnb1uiw4h+5jdKVUE7+2
mu5i8fuBtlntJDXPbzm9ZjeaXMblCPWYOGc8dPEzBIE39e6CJKGRguistKMJZ26Lr/V7oaegVQ2m
9wMANuW/eBC8hWlJqbKZmagLoIJcbPAF2kRWKElUbAvIgB/8SUKr+5kOsJ//NlArrGG+jRZOJzGQ
g9fLseeNJRkdLC2hg7/NA7H7qdnqaCmyG38FPCGe1jEkSAJabQbCo5kxpOzJ+fhM0+lTVS6BaRxT
2D+J4i4LARObfo5AhTLv6Rhk4jRZb9ueD3HgdNidm2Aa3jSHOQdyIiuwlah5oDzkICzMmDRRVWya
HAp3kvZ33GbnH3u2KZHFaVIzvOWu4sWoZh4wne2W+v9nIE4c8eeqZz151kLBbvA2bgF+yReiqaBG
BuPL3UTzM27lGB5o9zieykU6qlX2yOiB6GZ3DPwyz9JMUeMcRiFanlScpTDRdde9pp3STTs2cGZ3
A2iweeB5ZjboEfyJcyTE0zLVxRPHz6k+36WLaHdTSsoeGPDKSHUTru0L3Ru8gxPATLTCuY2Qs/IV
qi6FIBxiaWiSmavnxOiGfetzfqig6iEUXBlnP3HLTKQEiRv8PZcOLSJw3e17RQdXlqm3tjbQ4/BB
gXf+9O4L7LJ3PaF6y7QsJrtio9TQOBM0AuLRr1UAXRXmd9LzweNQvnAT7bAm+wSwne/jR+uOx71H
S5/+IzFism81cbR+Qw+F9+J0Xukyno68Iw7yhpsyXAFmmqnSNiZn050PdFWUQ6nuCfETId1lnPgy
otDnTTE3DtSO3hE082+z1ys7YqdjcaQa46TpJV3HkGC3kS+EW1yT4X4h2v/O/0R6kot+OlE+JIGW
0ZUoui38fojWsspBxXzot4kGPg4KUQNfQEQF/60WSgL0GEf+MVfR2+MAEgUIw5pjCWiJ48jwMkFE
p+LGAded7XCvBjqRJqkvRhsTe8NEXUPUa49tXlUnP/j5ewFqd7XVHqK9D1RbgkxkdBKmUVAuK19L
a1pr8VV85PSYrjYA+CEVc8q8odOF42aNuCVpjn9xDbaGharNyszqsJE/LtFWgKi371GdIWEiS/+7
vroRnCoRsIcxKlLaNt61Z72uJaGTGiDF+XrR6yRpFuFuci8BU8Iuu344GBG/McQTOKDYdprwAN5b
NAqKkDkH6jWFYeQtn2vWuBfMC5FtPY8hEQjrkNfvMsUb1eG0rm1gyFx4H63qNP7BxF/mnT7ZDLA7
du5jFBD3fv8ulOA35+hYePxU1b2FUFSsb4g6RV3gzM3mr9dH8wJuf06GLAU0uS0hZDRqx7xQRndv
M+CrYvoKbIQvIKErCUkgOa/N32mABagpIuhPb8wYY2XuBY6lwVka0RKIgTLzmhVIEvuaWDCj88no
9IS0P1hxGU76RYMqCurwmGDoBIeFwBxK0k5hbNrEW8k78aczmQjp9LziNCz+I8c6YBL4IR17g5zS
mmqN0OR+nkc6Iyny1MHhJC8ISDCNZHcUerHDh6IpL9vpBJBE+RbE9t7qIgNqYroqpIVmbkSQ407R
Zt8ogoOcB+uEvf/0+ZLTsM15Fd3jsv46p4q49dLFvOsiRHvh204XE0wfZWtwTfkr8lDH/fV/z50r
XggbKKtHdpiNtp0o2rajQC9s42QOq6Ej6BoVtGlPn4ZqMy72wp/Tmm0gS2vBW9SDi2jQXhJdRZBl
CoYl35SzzTCL+Ev81JHYnieTq65vo9hqon6PY58EnXdAateboRN4bCioRDcOJdeJbFEWA0erAQIo
KLk/ZOjb3M8UEdAorc////hq/7i4zK+ESbtb3xMSkPXXZDMtI88vU4g5KwmXEeKmXEF+Qk/xAqAo
SF4lLkjjqtJoyVKdtQjo83TWG0htusf1IJkUeE+IOur92/SbqvrB8Ttk2GoIFSiaFXXYEPJgBPSr
PhyKtOjCi6H1UR3X+uErC5aTvz7YhMa+hrE6at0utJCKSyMt5Iq5JtBbnwCEtS2/OcJTm+1w1bGO
eabk+QFlBnYf67NTWrEwvdn0wQAeJqPoGsUqkIOPFK3ZNfOtEtmc7bi0vfYlGl4ZlZwWqldbRHWG
ODT5xH1nh7f6/ArfsWNKpc2HpLbTt94TxK6FQxUArjBHyW96x4eg9PqvBxTgsCb8IQBK/6csDTjQ
xxcfHtR/xh6cTvHY5BHO5g2RXTylv6hH9XqkzvCBX2YSL91drWyV3RKZe1DwR0E+DFFFvkU7hf7c
uLvHf0ot3pJG0LTUEhjx+5RAUC2n2T4iXRKtkHp6d1StGBWmvrJqNWDDH7YJ+3E8P3o8zTSEgHZG
FbySzYIsWpUrfMGnsRnAX5OoBqG7L+C7s7IrULNSkSDoHXR1AzZnq0q2/hspJE4cqhYGgWVqrJRJ
7/4RvxaY3Pbvg1OnNbvECdawGlHhNFm5WasTPDNqtJA9inoyIIKxgwY8rUBRVctVztghsMMpv2oq
1+z1fqfGvhQxV/bqMxwXoTcSdZVdyHZFa75Q8WFlMWyVZXA9dv16PBeXs/5Z/7weQ9/DWY9hwOA/
yzbhXnwT51MPYSybjthfWVhTJKNFzoRsPQyU7E6x3T1Z5RJmOVhZmCyCXp7UDAgSget/UcYqSK5z
ZukFAJCXQltOPGKMGZQuFzcH8dV6EsyN9EnNyHy1llhacA/oqBgXFjUlUtv5hnsJwQ1b51AIatNc
n68lf02V/ykk1bi7WWAqPraTR5usdmpt0I8SMQsHqek+zVG8yFbVrpPXCwrVBmeD/gWPuXg8cOz1
Hjs+evO7ygTm8mfxLZWQT7PEW0SiaTmH/c8uOIrL10cDdZ0/mF0haVRwcDo4CVLP4IjLKSQI10qG
0Lcs8YpgpyXKztlzer4LmAz9xdVSgZnxl8C7Osoqc1K62Y7qNcuBBVj55uZkmZ7GvFPhB6xmw60l
RSBIYzEvAGvaELuapMzfrbWRnUmOze/4GEZTtZh13mLzHvv3c6Uy4QqJuX5PP6akYD3PLBE9taAq
BKWmqNYQPlrZFIcfL2iyW+36x97m0HN1CSIUOLjSlz1InZPWRUZvRkW1EipkQXZXgu0ZGTJxsxg9
sRoihIRNF7jUchWHiftCgAlnM8QG6J53IYCPco8C9mCF5Ggw18AXioLYNB56Fi7XunDduGtqreDD
62no3GurGmtqLPxIoYjMZx+/dUP4X2wr7s1aHYfxJ9Gmcyyfdtn5j9NBq0d7XNk5SXY/OjsYSR/z
4wIw74uVrvc4ZRbTebrikJoFNat9t9bFYYrMdsHXg+OqLY/z7bdGAdE8Y5l/i+Uxe/q6jUaFiQSl
ZDQKN2NCXbW6SlzH5VkHnhOnfhDQN8Bz4FUWnwK03IqWvmzndSBbQ1aD3QhMoJnM2jeLwFETJg1l
MD3CTqDU+JWdhupjq1VXm0xWiM1zg+WKLvZBpKhyBnL0LbWA5CmEdh0QXEyuuZE161HqovdCmG0j
pgcZJcm3K4jbqtEjdgYSPntvcLr54UIPTA9VxJUQ9wbwFvN63TbICjZFpJP0D6esesNxtAnk2qh8
mdIs5DR3MLpn2pcaQOr/T46FsmESXg3klWXEeNy9MBjcE8/A5Q1gsWMtrEEe09dNJsmO4mlxcjRE
IwBD9jl/kJmHnfp2KppscFCgiB89KkZJ00Mob1IuVhMMHvUkswMvNiHh6TOVLeDfOPQxrQkI5Mor
WEo0OnynLP3PyyS6PnNdsCTLLl4+CqEVlasn7hJ4cK88wrvOHFv3/v8P83V5E5i7od8y+vFJPRC4
CeweDh+caHQSBouBS1NIBHAWIco8BlLbatD7X3EQzR3QDoUDMDXt6hCDshlJsWD9E+ptGDYmh9Pf
x0myn3J4ozFdgSc0PqgQQ2vRs8neop1kN+1RXeOvWHVv2gW38ajufvCQZKz7tTovwDhAlIRRBgj4
QxzDfFWIuosw4ckFbqZblCjafYwK0WjMHicuQz+nZlrDu+mz+kMnHhj0FilEaKC/wi2I9Rmbm4dG
OObzZZ7It9sdDzhUDW/jiRgFld2x3bxZSfx9Nhc4k9uzIQWnwaHUqnI7AWOP5xC2mlWc0SHQ1MR+
fhZ3FC/54cH2/dN4dE+e3RcDu8XROPxRKXWuVc79Zlq9WthDqE+WxCSSQ4WRJSUlJl4fKGu+jB5u
7EMe7ww6RqqOQ8o0NPbmwfnRjm1y1gTL4WUXYysWbjJKOuHHvyB7WLFEscqTtVTfmeCx7EIJ0kYQ
BN/4o6B2pwTsUZsORtWvfdALxmXRN1eWgYWJe+5FqhtqdNcrwwGy9aRTiCXI2s5/2egiO7CmqsU/
P51GaVrxYifHda/26M7Fx3TF05mAYuqDbhZNJDLeM1goatIfgSdpRGT88idfDjnL3iWUYVSBmn0W
Jds6PYqsqmZ1Iz7pdbUrleOPKQSqChzAJcE8YFQQUZWyGMMzz+SjOor9KGmeiTTovAh+f7p+21hR
vRBuoeIuTCsrOmDivpMi5j7XNOxf+qCftL62x4VSOwqiYMU428fHhltwqX/eRDT0mVzTjlTSXIAn
hVlq/VZpbbEPdWPw4q63GFaSRQADYj5qhfrKOp3an3UKO9v+V06uk2cw0nh8DxpW0DuP4YmkpWL+
fg9Y6o1uK3/2DaFU5lo8fHCZha70L+xWm0oTszUCD4fTls6VdItWIOhj1+UvYW5+MjUPQZcL09IR
kQ4a3NJ6b1X6f5cuLW/LdCsuJ/MNsoGFAbzCaGNxtVe1ytyC0V1I45h/Mq7XZj04ZJTgYcrf+Kbu
7d0OpR31cFyZgjS99T0MREcqH9NzYVty7zM3cxscRZDxQYHzb57X+STtEXT8oxrUHEU82ETrdSs/
/yrhP8N56t5d4PnSzdWRnOBQGMjKFgeYzhd4wf27vK/uS1M0lT4rViaXTaU2lSNMDjya5P8Ow62a
MCKPF4YO7Ltg+Sdu69sE10l80GzfKpfX94VbjT0I8cu1HSXXhzzwTVhfrZxZDfgLoNLj44+TrJLU
nNFJu8sCBEKWHP9Rj4Qgx9yF4HcCFEk4b5W/Rvcn1wv/SsSXVBilt39vRt+G5HWbma4sEKZhrOSP
rilz9Pt9bB7X0D2d+T2B1PrIwxmhCprPB9kdWQKVPHvNtGfuecEopyErwML1EacVjfMQPHmV2jWt
qtxcsqsEe/rayPPZ48mVCiyU4dzDgDj98v1RZpXvlqZYdNL8kxsTw4uCGHOgeB8520SKGgzCQAzo
+rVKj8TwfZuuLrqmymNm5fH9WFe3v5izf606meUlmx2vhWToR9qSrZqUHRFqf2mu0uuWf90n4KBq
sKtdXDvKIGXNs4+vsKgezZXwpZEi+JRJe58cnQ9/w3KuRzwRt0NPTgdcIXfIuu8JzHX2T8BbiEVW
fnwWK3PH6hPeulXmjq3B/aAdNoXmmvaKEkW51LX8NlGQiWeHk7veAfS8TFbE/PvjzLCufa5LEvhF
fAyWPFaMdiOcAr/s783VhStXskKUjMtxX06lgfoXg+KWj3aPxFLBY3N7CDUi5r0eQ4y6BpzZ3COI
taNUHd/IUU68rzG7q0yUDVOF+Cz7MR7iZq2++8MB59ENJW1am0jZEDnQf/LOfp/sxebI6XzhIxG+
kvt6vjc74M36JIzv+/PckEzSGi3SQeRw6KpChptFPfzdQu4iobmgl5M5Len7zx0D/E8aNsQrs05n
2/IWULkfimAs717An45EyeqmgfKbRPkTcsXEZY6XZ2hnpoy7gCwG/B9xH5D/lBPdf6AezO+OYyYi
Vh85QHwENyqbI0Y/noA+YKjyGu5/zVGjD0SGpRjzMH+gfG2CkimOQGKAOo/6dHYRsf1043+H7vuR
Mj1AWOhvvfHalvAi+R0Wd3HLS3mQ/vf1aLjyfb6Q8buyHIRTq3qAx0O9MrlQtHBbFYSFcuBSKHrF
FDS9BvkblbXDMHv/MhLwSlRqlD58nTQAMYDDFibFzrEXuBPUR6vrF650drLRbDkhKNVnpQ7gpqkA
sZgj5N4a/rQeevCTnpsdcawc6hHfF3uPLEYM8AMrprWPdLVoqm8CIvaMBYk1m7+GUZywiL5T0wL9
NipwdxQ26E39F8KeU1eKvqX7KRr3O6S9XrkwHkWEArnHN25kHl3jYDGJ5lAIkX4JVLP+VFaSl0Fv
5yhn7zwawCtyuDta7ockXKJFb2lI6BoMRMlJWb+nqwqmlPBHEYf8SnQX2vri1g1hxvp7tE7fNKxk
8fLp7lVHxWknUcbig9+6evKa3Kw6q270jNNy4Nd4NIy6QKsNk5N+5/x5McM0Z9g5sgxjl9ePilZb
Ek26zG9fNc2sS1/O1ssBsXBGpygrKXyXDY5gs1DvJtbbkQOtDRQjVZtFQecprS86qamZhNQ1bJ5W
b0Mxbl541XtZfUK+4pW3LrhXuRSaUqL9/iP5TM0mK2R1EO2ATa4XPLbfWm9AyD43cM7Ko25dM0Rl
2bz9BUMHrTnlVmuYesO+4LvtgocYv+q28cGF23V+lY8yiUSbT4SVjSZR/A6k6uORLldZOHmWFm6U
lk6dMpv06oIiBhGUB+BcmuvcW5rOZDfnPJP3lIw7WiwhojXvh2ylpm57iJ8UuLZGnkHpv+8uOrso
0M5pY604NF3GiNZQHxynnFCor9qCNnwMQjt1e4f3/j+UpP/WaMwYGJ/6Abh4lTJKlr/n1o2rb6E3
iiG61/NljWiIaFZoZCFnASLNUbyCeGEosDAvim2wim+ZmqPdAa24BMLMMoshpJffKTaZ90BxSHMd
oiR4DBV9YTu8+69NpqRVJ9k94WP8o1ejSYV+JwqY8K+O2bAf/RDZ5RhKA9gZU7oWTkx1ut/tf8/H
d01DpdNPDgI7fF+YNOB7JcbP8EpwvD9gtrj3KpOzpIKXtRY7SqRuL8w6qfCEKl0OzA83//lo89fP
QAtFcj745qO4ULbRTTVOMgNCWzcPbeAQY9Rc7pvPEsvB5eDat1+hxzUM879XfbtU5ujculFF0MZK
7IBrCEetxQaCWnMEQnM8xLYz8nvNdHFebeBc5bn/geAE4nlCugMbDKdBHQCGqwCY2lC/OUj5mm/M
uN+qJlnsgzA6/U3WkfNrl9L+JYxCmdoBsNwIzCApNX1SARY6tIUpFv86+S6azGDJkdLRrmrd3nGh
M4RTZomMXjsJ0CH65VT+FUAWLb7vL1noZiNRRl2EX5DrkrKUUmywoSeHc1Nsk0+XAbwYwSDor6qL
E0wx4hQO55dLA31mWjbfBJcxVrUuU6mcJ3HWm4OCqUDEErlNAzvjA3xRc7mqo55+XfuxUxsKxvKI
fBIKMoI2lD3KKpB5rnjF/rjREVAaadFMw6AJ4EoaCUR/sqhSz0mEpls3dJ5/fb8asVRys0y72F26
opkK07mck8eZo+a4arwi2E6g4fGyOQaHbYnQlks9BhHSs7kNQ4btzwvLJkfROcDMMwsGEMHwQugg
ZYTTIGriY6T6qljV3pf37vDv0gF/bqD1vpQUtkVigqFWYpXYH2AAzHhTiCfdwOd2O2jY2Ej9sLXS
t0RAVbbRuEW6Q2f+biWt5+wvmTktDHhSgoERnyveXyDcxq1UaqqdnMQR2Of32kyZ3IikrMzKJyaF
MNfZC7mvLQcv5b1lfLxouhnkhJUGc9zz1KF9yTptfeBh6ZwFKC1hYxCuA46J01cw/apdmzf6IgLl
LBpgxIYb3mxJBtfd9cy17UZ/zumF00Uh4lfZ07f27Lxg611OJAIA/Af6CN9oKWGNva9H2wwROWiI
i4aRRMPSOF/M4iGo74I/hnd/xFuK1jZNtEpyLvBiWRoaTiqkNSVA+Mr6pi5v68wju/D15eclAAjG
UXL9AJ4/UMEguGTKHrw3K8mFXeNiHYpFkCqDd+ktW9k2/OSdwOemfZ2tjqDr3zoZeiVAY9ZAp7Ta
XPjZDlZP20oyEyqrLQZ3u9u0uhtuNKqGhYNwKv8lpCIbST7zEVr03LtS/X2Vh9NIhPLWEcGp6Ddn
W/WsN82K6/C7xxvvePqKXI2TmyUwVOoQMGpjP2KCbuHvSN4qK0c4EqpPE2+oRyT8y5vCj/opDSGJ
00p2CKzNROirJHGQtBl4iQdY4vQAor+gSgu98PxiK6wZ5hIU3w273Qklus23sIFl2jmeEdiSYHmS
Polsior02eorDtaKngmsFWDn+cnJK9f5cH9dDga1biws5qFLXi2mvWRUIAPqGKDJ+pCrMrwzZLor
mFhNsXIGSkSNri/IUuJ4QnK0HIqTxsTW3s77o4zcSrvKJN5P71u8XhCBg471RQq2dy0ICJ5gGvSd
TBaaMCOZHEWnbhKnYCAgiOYCkOJHETB2vBfJZCMqEYRd1H3ZNzbigvUP2uO0HYjk/0mfI+Pl3sTY
gzoj9bhzRY70ny8B7vWF7aYnevigc+mW7EX43NvNQMQQpffp7k6lFgrHLfXNdAJGh3n15LkIGWk1
zrSfx+GAj9ZdmYbO43ZL1rCkYc3c0RpUxpo3pOsHtcmnfrGRTzoxPTHS/oqR4Y8hfq+R0c3+nUvn
+3c8nZ1BfyFJ5/7UAsXJBdIRxhq9joOi4k7C98utuBby8cyo8lcOm54lumj2bBYMJXWRWD7wgPiM
H7/zklnVS6A6GR3E1PuqdvpkC1dD9npj7rHRUF/7B+hkCMgCxP6ChKwYfnA15GRLixMlpwH+epUZ
RM+wuKBuh5Jq43xhXuLnJBsezej38M2PWa16gSrK7e05LzK+u8N09XQcknV0vG+HSi23Op2xhRGS
YmtTHlSEb3lhnktEwhfsoVlAZL2XR1wyjMUCSOt0fSMrX4JDUSiNpyBALQuq54atIYo4CNzKHHrB
yeBGVlTCl7vy7HPVJf49vONj9AYvT2H6q990D5bwC29eSODEw65xSfPelfDSyHXq/+x0pgdWBH/l
EWtmI5kO5Ne9iRPL+0yh74LsUN81zW962UO8vxkmaTgPzPkybxGYm/CaMfUvBb6x7q1I0LADhruy
3+n4USX1iubXY1gME5u6R0udANGU/adYCzmmQ+PTJcDrMtrCPypBnyszuBblKsslw1ICNqySKTME
UkqmvhST3qDEdHfTw+Q4Zb+Wfo/eRu7lXd3fOqnOdvVJ8jalK2feA3tqUzQb8DcWyjn3pAi5FEnZ
H8HYeOD+z/aZ28IwwYXoo60kWgCUgjTcOArkcpgA/dcLrwx5IByLEGgSnx9hzwykYdViWQy4gf+O
tlXWJEDcH5jky5S7T/ui8OLSwkrEM9oNIm7dRADzobZtM6kj2pPwKj3hD+gZ4OqZGTv5HG1coeOr
9HWmpARRCSwBWwQaKHRufxl1TaOwhzwTQhb4jrDJQ2pdox/vNixjBzkzrEinzyvEodBNsF5yoRab
sO4ADj8hdSoMeEyR2jAs6Ves5fa7t0FPVZFKzeQa8ObfR/ucCjJAE8LYQuZap6Py7JHqJltfio6C
DlXc2X6cv32rGaW/g8Ue5bUSP4y2ceGz4Cvbzve23kbLSPJV7HAyh7MHYP4fPa9nrg6afjVh/lgT
XyOHY2qJ5+Vdo1nySsJuVj+NZWRpVU9+wcewR1PYUxjsshIoUcgUju7jqgCBPCrFu1CeSag6pQEi
lfnT9NRIh+jDEyR3Jlikre8LHviSicfQB37fBm75B0yVrByXLcxa+H0nHjEAmuxNKSfHYqcL0NSI
pp9p0XzpOfZHUoysqLv/daAaFNaokWgRkpegv77YQx/s+UsXcPycrO4RcS3Kf+LnjUb31ysQWe7V
vhv8rI6uYMYHtDAPtEvGD2SYVjo0k1CJ6KHFDzGWun3zmEixN11HMuqL5eVwytFgwDmXz7P+JvI4
nRJF94G5xXPzVg57mjXwyQX+vMsgW0495N37mN5GFrB76fcUKCSUimXs+GyXnBG7v7ANN2/jFIPG
MIZwwyG5pH6n0Z38ahI5e/Kscx1EOhbM27q8g8oAN602jLHiTdjqNsOa1AenUshOegD4byRbtjhR
X8WOGGMYj0ZZ4aQBA21K+5bewDC0QkHrPcPqvvZV9vSXJuJD6k/P+JrLHmHHZM0Z9n2iMRo4prjg
g3kX0ILyt6uGCwQPeFr+v+hQZAdgMR7HoH0ZwQoP89vu2KpNvKVMN78fNLTyF8EekGRs+7wsLffq
D7wlY0xg0MDS3eRpswBZGpQ70JCC4rOA0PDq4/2AFrGkdWQL1Jrq4N7Gije1k5yr9uUXUH1A8Gft
BcOYHHnBXu4ULAOaR3z0MMZI2K5UJXB56atmsrkHE6rDWmPNi1chhEKa36FEtp2U2wyVnTqz7mf4
/CWkHGUcbGGrZRQ9p41PfiFMa+77ouGYlcORaRMJRvmAksVkv8/eX97J0AvsMUtoJt6N8hbZdfvO
LIDABp/m5ZO+QV9x4DKjDzx32xJOTqn0B7JJm9Tg5+gvMVfGyKUs/O9L2Xg4OoOH3JpzGpWmydJ4
Y8E+mVYHXoO/kjR7B8fEJV6928fn7giDakkctJmQJcyqPyAdrvpUUMnn8SusTO1gxg3UWdZiJ4PW
wzYdeddv/AQE/PszsnBIVuE9ffeST9/bmEg1A845T3AJFYMW77Vq+7r8akY/TnoPeu8dTAsgqxy9
Wal4AnIO2vB2X/u1YiDDvOESAjg6BkpIO7nhJnS6YGoSF4h1fE7tgLqY9Hj0FkhVkN6dJKrkT5L1
3j6/oqd+JbOW6pqF1jNTxUyQhpI0D2wB2hwodQO4E78diXyWCr4vv5MLuk680ODh3hOENX2Dqa4Q
U/+NMYzrh90mRD/LFVc1+mHtZMLfuDyeBreAZME0/eVdkv2IeKlibH0WsmBO89IssL+g81fw83XM
FAL06XfWEFDV3wR3hmqKm9CixDiLJ+j2Wi45PkDQHXO75pP9LRhK0gT9UcEZuWeemJFLOmqh/xcs
yGP3F62aAYAyMZlZHZfOB9EUwEeBkmmVWCTkGlrVBwSSY3J96JFWXcTRHz4ij7ce0tsbhCM35JQm
3uWyqxbjWBOOt+e0iQCTNtjyoPRLu5kJmQNk1tqt+sCZaLk0nuMZknXm4GEW0FBD1oX9Bcpc485F
HKcLU9fBNGu0bAJByxbX9OFQKKIoLiDSa5YYISgROXUngyOnMgcrufNnzX4e+rxZYoz6jMXXYwuc
klWhvGFnvF6h0f6IfO010qCfmxVLmr5ojcx5wyqVKXLrF9MfalzZi45+RpkPS7b8xXo3CxJ2G2O7
7Z7Ma0UFT6rOgUSoZ152NHBbpt1ZJuC0+fEXibSST1hSciXlkNPgoKOwxfp9OOWLJ5G6tTZZCx5e
C9H+jPdti9zoXYRwnscTSqVe9It6QVig9I72ft69ZjrX+MLwFmZ08cg6OnWxNZUGkkdyzhUwXMCm
lcFLz/MapNl+QXMkDnBpYveoMUnrBeXrcK83eEZFRFJsDAOXVe2dUBvaFX9Y2i46gl4fdpkLsszD
hV+Dpbg1qSx76yPd96MWL21X4UZFhDOE+udAeomfYPhIxm4KbAJJTSU4RfsZEkutgeEI/2YZzbAV
bkFOLNkLEH+B82M3CLHjRLJGv+UnvP+2GhpNdEsvc690neW4kaMmRLKgKUtjCzT2zShA4AxMdxpP
YP1b1aQQj9tyYX+GUqUpPtltwexIKhnxzbg1gVLoXnVtLAFnTtoQfERAqC6/wR5ia0Uqyq4Swtm8
vBSX1g+A+7jjqCmvBodcmnNrOr8S6o2ZxZQa4CfbW4zJqaX/L3rUlLKneIKHzAaPjWY02tpH2hbb
IAoauHbZ9fKbXzchyQMd6QlNv2gKE4vrvANenODtGHQPsrwRixhz6vnD1EtPOxGDVkLrjRlNzBc4
3B87wotavFZvfBrJM3cxlB5JmbyRaVTnrDz5VEngFL0vcZakKrt3mnOcqWGKkPA2nW/am8e9GDYZ
at+Gy1aeGPYiCrn8okb9jFxOQrzhDwT+Psn354I9VxgMeIkogHt866moFWZv5WDtCItUw/IFTpek
SFd/t46/q0rcGANYCquT1SxIR3lqjo7B0cO84ueYGCG9FhRN5BbwYUkBR0OZvJYRCwElxephuRRb
LRwekZj4u6omoSU757wpCiKuUvlMEjwYkqLT9wSQ9tzYk0Faubh/a5DMKcuaN0oPj9+Xd+GTnn3p
+B6CSCcQzsbgR54jU7l39PhcqoabvP8y5JhF9ee0pIAfFT8RVbft49Fe25olieI6S/J2D31y+LWI
WiA4bgfpZZbR2hhGJPK6hmfv5J0EUJVjdNaCPR0QS6u/NgMWSZOrfeV70cCKR4h9Ifoos2i82RI5
Cv5HfY8oqJMNdPARiCv6viMofmQkmxAa35L3KmJ+4C9jBXfHTEWhHwF/l4PPO1Pd4zAI3Z07Km/4
G4IIzGt4seJADDstjHKxb/4lJwxj+VrDm+mNJ50VNSJ6NfJPNMH1yp9av+9lLNAFBtYONR5leDON
Dn+wpTmwdxzcL3oK3zwW5jMxTxCDC3Lu3dqg1UiRxa0G83DgqjrVEWvaX7E9b8VnpDwm5f115QAB
vFhOth2qejA0QijWfcnZafot3WsYbhQ+3O84Uv6BB1IOz697KP3zWWW1VlLY0C/Jnu1mOh8I78Md
Yjxz3p3trsM/2c3RNVvkJxcN8aFvHDNdRhUMQuZ+ICocqOQOHW4wOx71DzrmHfmcWdfY6bYjV8KD
frRhvvcFSlMPUVHtYTPLV+aEtT5Dj1zFLiu7Yii7goT3u14N3dBJUKhNFVekkjsgceC0qrGrdFtP
ikysdq6LR7HZiOAyA27AFU4l9JNzQ6gMG0kGUfyDdi8hR+D5MDv1VEuN/99wZAmy4OxE3mACeMnZ
tFW1qe75MWoadJUfU2W1dxNGy/jxStWvpRvnYMJnbktjAK7Zmi75jXZQgv3J4Pu5pwkgeRA4Yb9H
wjTiz8a34p3jLUaqX190mEYtYc0OkbZ7xpf908ShWykx04bVVzF9WPUckfLZIbIxa07u445QtmW4
1yUgHQIZHB1ybyQzGgZN+38/gp2DFx6stxTmLNlqbxeWyY6NPNeU8aGcB1z31E/VM8TpNtRlVktt
smW0/CCV0XItPpAz6YrIK4p7j2BxHam7msVGkpn+tqN+dX3eB8Z1tEVE4Omxq8z9IMwF1OOpL7lT
14smuaJxJnxSSUh/oOZdl9Ks6m9+xErKrYA8fhoZMZnkMchN1d4nO15Sp+IjGLXbymJKnTzCZXsn
B5T4UbuQvVU97D+xsHnTem+93L8PLf/2Z/HcysPtvcI1+948rvpGwEfen9hcg9zAOMcB+o3+N0do
c/H8xOaNlF2PZiA87UVYcrSHgkuuxp4jac9evGBXg1dEHBCKxUvNrIGd5oip2BBjjxbnGXuqn+Uy
WtZtBXWkXI1U0pYVxFS4tRnaw81fii4fWlc78XxwbIBCbpSZGVZX2iKJC9TMPLsabWi3lbXLJ20X
FLT5ZBCQiwtrvFTAQL69xhStwiZkEOefdzRJzTp1U12lGKZMKowSdxDENcGRJ5RENK5n7RXvso8c
F3yYJv62vh6phPVD0CrM92hKb8/KuByXBrbwfNh0FQnAjB2MHyClSaO/NZO18VSV11+bS/P1kAGk
hNqIp/uaf/kNJ1o8nuwic5nvACQJs/N988qIHA2rZyckJcLxFTFRBXZnRG6ZjiLl1ZrCqIyqWXQK
B6gAPai1H7npc8Edp87a4+FlJ03Vk6LG+0/SvG7FPW60QY2Avi0ADSBino61Z6kWIWvLAWbFonTG
kd+GlW/ZFLIIkH6afYxsAC95fvi3V/sy3hWeGU7DAo76tYQfOJ3oiWtPWuNiC6WP7J9Z1fdMCkgJ
+Dg9l0tYkN3nMBcs/fJsPO2Jcssqhf3OZ0btK44OkrAO+bwbW8rtVdcW7Gbdco8F+AD02w2JSh7X
oSl7tjxjehnN8RjdpYaOyw2g/l3XiFu8h5YgGBkxvuAQD80PVafvUetVPM02BYOjNb9EfOj1Tdg9
eWTrL48D1cspXcziI3xdBt4AgKqkBxTdD015O1Ryfxil3dCgYJXrZ/FsMLvxg31QJ5hhZFa9jWsG
dZY815FZfYtJYJ6sR+6UqbkhSIhZUvp6JHRBBLMTj74QPUg/MjuVdkXerdzpmBa9TZ1E9RVgoElR
RFoSU/keTGBdK/6v4oCqzR0AxVJfqDEAkCHg0jmx3QrxiA/7gQdXkGnyYwXfCnDitPl9W8lRDGNq
3DBNhmsPSk6LiR9+puXd+NaTyqWIZLcoPVQy96HWj3cWsH6xd/trs6PH2Bl3Q8uZXIvuyeB1EJD/
om9lDvbkoqRSSj+ttOYt+qOW5Qm2SjcsG+TkXWDzKqIJkIdLGP1WwKS9yLyRfBZNfUpCUeOYZNIS
w9ASG1p3xzgAqXWsDa5f9cdHGDTnzZH/J/tdUMCphhlVUkPEFO2iLDsG+qvWYl1T9tiQWvA2MGX6
q8CuAzSWrBh7lWYhF06U9ic9mmrAQL+BHCFbH99vPrQ4Y2XgdlwZOB12hL7tqCnXYBYGio76X0MH
mTtBKdnv4NjesdSkQqgBvWRpPN5a141dhZGE3QodLY4EXflHMm/XcY6AwC09LcfWsLyE0+XYfYvN
Rx9t35PUVavBIULrPUoa6LfvjTe6PUjCNgVidfPOLN/CSvP4dXLBMNaPnw/p1vS7F+9hm6Buq0ME
BuSHIUJViPBB3R84uhBmazPLcAYqNtuWJgd0dysoC3x7yqIVTXx0ztM1QDgmCVjLe8CIZTK9mlOU
nqtX1M4iFQhOT4Fnd5uvzrbaZEhrOrBHogdGsiRvBgWZCG7iMtfXagGRohAaZahuPuasxifrUoxQ
CURdd4l0DycGp5D/CISwKqNpmg3WalbFbT1q3IB2mr4s4V8lWf4WpfxJ5ZWDzaWSFp/sZ4futA1I
upb04diVLt2pB/zgYiM5VSTpMJAi6YDQ0EbOTKhdtCBKVUGW/A1QK6PoI/Q1Jw/XeKsHGMAD6YiQ
zPnilAiFReUjSjhlQnL/T2pBNxobLIwCsr0E52KPHpcJJlyVSxOcA0eflSPB8KpLqAto6pv9ZL7j
TFVxQ8cB0/xm1W4AwwScsIxf+w6uZkEc2xlPMG9xTdaYKIVOigNNxMnhCzVjv5DU2oq/pZsEC+4F
rgmtXSketrnL21tkpdKuKgue9dEkJeH38gNPQ9x8AezkZ98uXPPJwAu6T6F1jzvUlKilBc38+Jko
YPrSjgb+kmJnS25dRhnZKsj1es5NshQU/huAwQ+aesjPMPb3V1PNB+bi7tOKGRw5+Wbl05OcHu7r
Nqua0PkaIofI+hYXUWMc8es5QxPK6BUkSv94/Eu2zIGqjrNXdQBO6UrfggSX7VqFW4K//H3vYWQT
Q+TQEPwmYU7G35e8hJf1mFvCFYoKAxlxwjGUwhF8Qyn5XANoCk/LaAhdnhlhDZIuVeEY7vsRt/pr
VIcYQHjgNFNVeKa5y15cOSTfqeprUWgaI3X59GilNgewpsVyO91D0wcL/Vl/eZCrP/Z2HJBMFhDx
5TYZh3w7rsqxuxlOXvVs6XV/J1u0m5OTQF7Q7+2/bPgzbUAR/cRseJ3Znxp1fadsfTNWX5HMi+/7
YfFBDehdxIwu2TipMbqs4Ia9gjvHBDcki/PAHpOfDGXt9e3Jw+tiRzrF8x8xWmqipF1C4ERKIlsR
ybd76WbSmYoIa4hhNDMx3QVJk5vuuPba/wC/+HPDF7vMTgQvpyR5oqVGke5vvaZE/rzCgVAbFDtx
mDNeD6+oJR73au+HL2/vGY1Py6JtgwMnFBMFyANbwC5qN/6QDSnqMUD3hTI+3o7VJbIBStEinhNP
mWdvUGByTCyYzv8H6DoQ4rzFKuXAiIZERirJ+Mrt7jwathFtaTwrleBDPeCWuz8G6z2IzXdt0F4D
Yj/rBywF0nSyDnqu0GMnfs9ogkdmplpFVQprasXYJZCKeJ1XPr1xq6fX+dlLCRUQhHpelkG7NnCg
YzMLdP1Oc34EHWfxNIOoZ5CanHH3ftMyeTpxcpA08fzl+hXpCocW7B877NEt1k1WJEIMK1YwQAeE
agBZeI+afd4rJe7ga/F77pug3xVarVNcyNbUNPPE6+ZgvanYmtt0ZAOJOKGg1tQQPLDzpZc3NQfk
7BsnTsBo3PbW2LWvnOJHoNdi4hd/XVPaVE1rNMXoRJGxDOdeLmsjJYU6gtCyH+0X81yqatIDHOw2
28nARC68NURKI9kTIn4Q1HLvrwrgjbERkqUYglpIdQw2WY0MZ9VURWglcXP3ELIq1kQx5Vp0pbzX
wpsgLbAMXnc49k0SDu9UwH1ylMOIVK8Bsw7Jkw8HIZlSuU4rwyQdqG69uvLVxSCwWAtn1u76PDVG
xZYWnJa4pyghoAmbZ8dHAmF+1uh1TSOFRBJn7IH15/5qVvH+ZFogxgq0j1MdpCFoZiTMb4df44bK
W5VhjYO3UiDEO/r376DzXyq/AzXC4+M+rEpFIbUeVDsj7E6Ffm4ekbaZV2B074DVAmclKEKhftEo
KCGRwK71YrrBxqM7vn5zq+WFFUnUZJ9OuGylro3h954f+VV9qn8/fsf1MMBFcNnjebYHjftDuBQT
SFDLXHJME+EaXVJP7PdnSiQjpoTdG6/56gpOVTK5Z/D50iEoQvnhJmrTtHC5AVCDGuFr/lAMEksz
ioDo4jWaS5PfJNqYUL/PYfhEZGhpSjeFQYiN7ALPImmTv79vatkCE3Zw1j/OAZdJ4jhqI3M2E0lt
0xsMBNfJO5ex+f7jGX2i18olsfRBRSHDBqutPoMkkzclT/GtzV5fcrn8WAgyShn4o0zJfnr6k1T1
7RB//rWCs9fP1rTuKU86VrRAGbsNOm2PvX373QIKL9SL6AP4xcfk0y4fLp9wsz+4m6KOOLnzQxCW
vZ3E4qclQp3cpiZhNJcIzEcbHvzn6/25YanG9XmqiWpxaCfqeFxEpjjO5Y+ENG5drkKc4C2SSXIZ
ztL8ajXLPyobUV1+uQAopBc1SLeA/ae60sdQZen3tlcepCVdEqAK1v45v5ZDiiDIRYAxZGHbf+KQ
pgVOnprwVop2PktcAv9ddJGBltnaFhKKkLNyLmhT1E7Hd+/taOAFRhHxU0Cw/3b1OfTT/y/iCsNC
xICWvSrCEofCwA3yJUY+pBTAR4CD11WI/djuA78h4G/9uvDZQyvcCetx8crilq+6L0p1ZyJV6OtN
BVGWXCD2pyAm8ReOZbN/X7v0QnFTmwQydAo4V/135xtAxkJzK2cPeFPIyIsnaadOXmaKzUuxK5LH
ymDs+xVBWZk1uYTI0h5AzuQpzfJQR7Kn/PxGMXnhrFdWvPmv7fUz6pN3od4VhaRuwx+niz4/BHo/
Eru1c3snOW6wbcaZyvm+ZX2f26ZJIXw/XiTEgbxj4o3ePZ0SL36NASf2dazhoqBK/e/b1XWfHRrF
e4V+G59rXJgOGN72gi62ETc1aKEcyepD7SUzJDL+2kz45puwxGIJFXANzn8MXpqlcxubTV57DhSp
MDFuVYJReQopYRtYIceK6GrVApE1Nm14Z05rpxwp21Yy7AubiWeES9zJnXKTyNzjiaNGi52oAtIB
7cwfotB6Qja/Fg1+Q8teeWjs0uwLkMrn0GgcoibwCwv1LOCe0SxwDp51bZ6jkW8hxLW0urL1Ffh0
Lod2PDeAiFsx02ADWOzbi3UYUN/HPtaWgMDCWStqB6FtVOjgnSwoEAb2caW+ycYqpFVGGTfp1KB2
UZoD/MLAWKpvlzC2XoH/oBxA61WHc5nHIAjcUYv5rReRt6W7XI0CNTxy6p5vX7ZdAwdrwnUZ+3bV
LFNIyXiPhUt0OdZdKbP6Tm1sJL+FAjGL6Ornl2Dd9vcjtaC87CwR0e2jmISoOeXkx5fn1GEK4J2S
HfAylO5ilIcyJq7TGa+YEERrtvZU82kSAp9JMc8aHtJY6SCRpZ8r2iHHiT7uraZk7xcBNMKNlB16
gEtV764YOH7Zkny4DVKw5VVbob4k9pWxKxnEibXzWcfMwg7ruzUR8NoNCdcIeZru4dWWZhBWG8pp
5PNQUSZOZTiC3pYcEPAdJuj1OMXg7sRnh1nfZYvhRlOAXRw+3sqpOPuRMhPEpmxpofRZasi8y0sj
2HxdO1k5X2XHqykui/E5NmqapUh7WHJwi6eUVotqt2MtyY6BSHqx5/x6qwVUOaTgmqpvh6ITdQ47
Eju/JB5pKuwO1U+kIabGcg5+uk/W5ynwR6GQNkYR/ipVtpL/nlibe2ONqsBDAfp2JOCOJpi7RVi7
JmV0xjxSERXrnGC3O16n7vTekokKb+AwiPP+0U+dt+fE8BnfxFW2seqyjQ69v4NSdJhCSErF26el
U6uAlxT7pyrm+QpkIOUhjoOVmukT4PdQ8SEaIwDv0HNtcOHUH6tybtzYSSh5FdB6bBtqshsEH8Ph
pNedB/l2q4YDoeywK4Z0pKhRwN0LMxECkRK4j4EGeKuEYGikplZ1Pr0lljpsrkYe9FJ6kKDvHoj7
CwRIl/IQGLzZ8ckWfjuEsjgh+yQE7vPZi76EGtyN/BfZYvji/avpeMHZ8/V7G/yCitzJKKSRCn1D
f2w+kCye8Xa7WoJlYi683vW8WUVW4hivlshDlK2f/FD0aDFhFnHemGA9ZT60ZFACYfRJL9ikNa1N
EQUFcd6thpXeIQU/4GpK+Ndty73bVKEgy6QJIrlaMR24GVhZ/Gfe6i6bXRXwhnZyne1MUl9fbmuf
4dlLo9N+9Ph4UAtzWZ/MJ2XyvPLNrBkvLSV/rz9+P65Fg0QX+9I1qmXEs/qy0TfoWuDbPdw3gxgc
yy4e6/wXFsYeNyRphvoD73jpnNpNZhzGNrhQG2xrhrDtct1z7+ankuiRvMAiD3ZVmenQ1GcIGGBq
x2TdHfysDrfESoFu6cCKUoWs6Z2O9UBbrKREJSkrqgFL60w9ikke1EaRxA7B6xKBnf29f7aIdk2v
dyyi7h4Bu00BN+g/g0+b++RA687s/tCIoZFMY/kbVeVI8PZrkI3YaNPRiiheRuLSPWsySFBx45HV
OE8yqwN7ccSDciWQYehjfr6p4M+0Gen1btUymhK5QGZ4NG3go2TckxnLh4iOIHnBsmQiWKBWmyQA
pTBHWY5mQytT5RiEnxUx5KQ/gO+hssRGPz2FxihSnwSafue13TOrF7OyrOFO4L1xZCJiYXLAlrzN
NFyMlLONvZ3Ck6vKIry+WPzjcZvWO4wwYeJtI9LkQil0BlaV9rR5xYbjHFII/Hc2edY7GPUSRfy0
LliLyF2z+yufixm/5PBVWOc6HGbyIJ76vOYk1htmXe/gO1vUAjBuzg/M+MPjHjGiK8XFj5sZwN5l
SJEqZnkYy9FUSH0WteMsuL2Mfl5sVFi2n0cwQQhA3QFzEFQA1yT5hHKpUCnFQgzd9U9GjtcjmfU7
plmQywudGTpAR1McfKS9lJpi+LRSnDPVJH/OEqnZ/79rhpY9w3AwPcX/MuKbI0Dn32rNYDMl+o1I
MRl+wLtM3Q9NXyG5LYgB3LcNy1f1V4GIzetp1AsaBXKFHtl81DmhcQWbOiHz3xvrv4mXLe3uLXL2
ANsabHk607jXpGxdr2YJCDzh2mkfTeAPh/F/iajfSasVOtBisOGV7Vbkt7Z4ujc8NWMiAdgxpbCz
gChuWs7sD4bwWnB0fEnjmTLXc7MOguIe0KtyogA/nlkHPYQq5hICDBIXLekvDvH7YjMeM4BPBkEu
1uAZ4iXJxOH0zwcC7ChTVInA0ujyycZG8I2Ysq1DCYK6rcObLcN1BrkWkbH1GjFh6kkX+O8kaAnc
FmuznM2v7Nc1cx07EKphbPTc4rBSiLDiAu1JqffpVqbY3GFdqrfaQO4ZukDDt+Wjj3GSncZnoaK7
QaGLM+QOtrklFw4jHRWQew6gytByrf4wv3kxvSzzyJLD8F/pCqHGMiGgQdk2NMu+0EaKIcuoXydA
2Qzy8ZA7DgdZNF7w4zwrNAy7v1cbbbv2fPqRFjUzcO5rFcJz5wtvV/fSmon8htHMFeIA6C3s037f
nl9PXp8338hatd5+x1XWRwyj/1uf8v+LgNpa5bDO4mA6E5TPR69ZgZyUGYZXLghSSQt8ADjmDTAu
+Cpqwr9/rKX53gKzEh3+VNE+aVVt3XV45okqbGUbcWeh5zGNdIH0oU8mJCbmuf0fsal/o7eesGTx
j92/MyzWzHU5qvvRTbXnIC+mSf9Th9bEWO02QCZ4wWSvC+eyIPJfasz1phcqtTqWpDxcOXr/Io15
DgCRw1UlEiYXXkTxOEhU8NPRx39Hw3v0dPT2Tc99CHqN05l58NtGcaxPsS6Dn1BdqOyOEKoAs7h3
K7XY48RP5Mf1SkNLbjCCs3JmZhAdlnopiKvlEuFc5npqcUPtfvneNJ4r/8vbJNc3PU/pKD/m2Gke
sJsJp4o+ausDD08fWlMALtucGDAUcLPgOD5WL2PRzBQC0t2t+Szvx7VqYisJ+KPAoeX6qub7QU5A
oDSnGYe2NnmYF9I8he/rj970fQj4qPNp2peyEAEEuhDuQ2CyeGvdEWOv6lfydJF+d+sVxivN604G
8OZtfeq8lllGfNl7sacdqDDBGwOmnk+0BqGXvH0v+NDakau4vGcSdsJMpIr30omv2XJYVmtmn7iJ
0Gni/t/aIa6yC7OjZGTjXzt62cB9BFj67LyyBDeEq557faJUzUxRO9ZKADWsDvgU/D/iEJ1kZ4FD
41rY5b5mG7Nt0qUiz10vErV0lrj4eqdTiDiIg/LsyzdyMZ4FCzQ+9yyviCG778XnB8gOlg0w00cX
z/3sjj9XJhczpOgi2Hz1NeSOrbgy+MbDICA47PJSqpP09J5D1UKDncxNI83xBd18CjMqOE/PuCE1
gDwuqQAFqUAPZzJ8S3EFieyuiLKYgkRq46aAJbb5KOW2Y2QjhlRGvzyA5UVklOTpJpVR0lh8/tRU
QvXfy/aQXukKh+fotkNT3/MuUJOp5+OYQuF1H5eowZTg0AdgCi9b3ID7XTDW4inB20dIZQ7j8xfX
5sveducvwJ9ecxUOyDhV9FM+xWzdhSBL340UQmEWa10mGYsTxPlWo81Fkpl5on3lYNbrxVX+aX+O
Y+iDzXtDKGKhC5kOd2P5vslMD2kgF3gkzpg4SEcgQSmjbUBHc7HvHG5Myw/GAVlKuvgMCMxKkN6M
RT2qDM8o0jGslfxNECIOTQZz+7bN0m33NEt9uimfn+pc65cDKGPi809XczPeA92/bjJ7EPJ/I9FH
soj7Gz+f5ro9/LLj6VEHLhpjkM7x1/DMi13JSiB63ruwGkUc2l9DytmtjisaSFdFrsXbdzpOnLdF
2L5YijQCmJ0PcMxi7a/LDXC71JkJ7CBfaRAKAH1S8f5ZXklK2kyTQ/Bx/UxbeiSJGMu5zLJSl7SF
S3JhBeuOXOH5kWbgXko8GGLCOcVtIJh582OLjg0LQsLF5kHJ1rl5//neXkvMZIoNJNmctAQ32u5q
pH2Jk80Sx7aJM3zkRlskjl6hRtZCeuXwjXU7KCKXSg+xbd+WUiaaCZxO1iWAYZ4oQSTYItIN1OQ0
xd5UoRJKrHnEgERGcCVq/Tm9J1PHkVMelr5iNpVEx+8sd9nbQJZ8JoD6CX9kXw5PJdygntNw1Gdh
WMBcC+yevlRQv9pBor+0heSG+pQW5Z3Tmugc5NjYEd6xsmW3yW78IV6CxmmlGne3GdIfe3twyT1x
HXUbiFbm8G0PP2oI2dJNjyl76pOj2eyYkGPbXLv1BGtoHXBYRcKt7Gn3eatRsnAWMoErYeE87yBw
Au5QBapZYpf5ROheufKeoTSJoQ1uky5zGI2kBb8NIUbepiUxD1VvCC++9C6XbAP4JzYjbjINlv8Q
cBRwdnJxcrf06n/BNUhMSApWDeupLhVIDu6tuOI+8snCgGwsuXQQ3ANdAN5hWY0GgOsybnhMrVm3
LDNDTR8vjHUV9J4rQUKcx78IU6jF3vPBC2rD633nVREoutTU0LtIg65onGQqzrlHj0DiH9BqmHaD
vni3eLqjGWlBbnajSCwu/mH78wkVavjooVtTBHIxTSz3GBrAErooR8H4KBP9i1pWYDzLAGoCrqEB
gTwi61wcGFI9WIDV8gjac2R0017BDS/Wogt7bOJKF1bhWd4TET+nO/U1ZmqlE/yDACSkkNXE3Clg
L42WHmkjWU2Na7WOLd7w9Hogk/ZgpatiNjiwgGfM9zCNYZlTpYluZLlFn6ElnDTRb+I01AZ1snKX
B+WRjFYdR9MCs4RzgpnMH2hmfFkqTYllMLEC4w02wdknSg8ns1ec5ZPIQZybOvm3SN8ws2URc5lX
NpP5BD+fdYaxYORK+sCaunzpV+kP3ftkGlPcmMbUcwWBJdj52cTGjSVjwAxEdfUdoFRTgEe2oOjT
n618fEOWZDOEY91+ps37ojhLpT/giUoZQj3AgDfB6ehjSgFSJmDlR4YCnllmBqMsEA7MB+G83QoU
9DK/54TxTmO+p1d6FsH5k3Ug3ZbHMuupG7eIuoQ8IRkUvLcuy/6aUTows22jtHiRgw1zDQqaXlsH
BVOtzmOmWP5GoUlX0JTuD+pE7/e0m77S2vndM+lwBtJxhb78yhCMcn/vk5EIKHT0+BCkOefiXctc
ajin2HVkFJpHqFMJVoer1KQ/5uaStktBJn4TtWCZ63mTSS5wu68fyX9LfKHPxdVy9DX2H3Rmi2t1
tlwrxQTQPmCo+0pqISF6LqtCy3euwulupzIg4qDfcnmzRdTleF/2Hxkvb0p+RNHw67X6F8OWQjpJ
BFeXr1xUwEmuGv6s1+f/l4Fi670CowexxesHdJmGmDw2ws2PLHHO0KfAbYrEn77lkF8iM8Mlzv0M
4w7K0+gI1Dny5ORT3nK2md5TVYvwOB6GxETb1O/mMvZqpa+XRdFteZHJImh/skJzjYymiRGMlgCg
rvsmvtoYjFdshY6S4zCqfscalAs9vygD66u1B1ixQFwZQmEAJVhSWuGduN2vPwU5Ejs6Ci9neANC
somwukqP0tAD5r8fGkc5wOCCkTG+rl2SuNmbIt0DNDcBMz3Ix8WcAbYJ90soNjlbe92LSJZGqH9t
UQWeWKj/AO753yWBQHU9F8yaJW1pfH7CMBXQ3sXyfuJorS/MAnQnioZqrDDgf4/5yKGQDau4ZfbJ
mma0Vnbx5htAVp8V/eQLQs5PEVsx36SSOaHYNH1+b7QP/bthVqO01/nOrxlDUbrgMhuMYxzsVyYW
ppGA/icntFFIpV5LOczbEdlC1J10aXOj9MOz0eIs+/+EozqyBl89PTL7/30yeNq7BdqmLEvKxXEJ
qZGA6GaMRjr2UF50MWWwbQ5/PeY9xYMaRE/K27vF4HL5lFzFyMoZlEhHfGNaqhclF3JvBzEJpya/
bR/oiKvBaZVwuHzZ8mH6n95oSgHq04rndv15vCgSRCYCT88m0xFvKTFLt5jcAaD39+4c2c9enOrK
+WWIAy/udfYLP36iRtNk6Gbuwmc3pAMJyqlqi38HZekTxwrm7AZ16jRz4J9KuzxG7PGEWkwTBulO
3rWSDLo02Is/V8V/wotbOcAv2cgkk9G3/19apsumJ67hc23K+rADCkwbWFUWUR1PduZ1WhM8pBjh
Dde9LOJgPvX5ZY72vzE7hI+a9Okj/hCROsX++Hdkv3IiULoAXs6KaXSKEdjWh0PrlCXszZ1W+lL8
CzGE8nfbKoROPqNJEfR/I6UyiKWhFaYt5cVwbhR45/gpWNXipE9AVJsLkgU2bM/07czxNICYx/99
p9jZcp++Pp93krY/vYYqHLFSqD/REHPCvGqWrNW03qqOHS7w0q5d+5uibc5T3JcInvN5YTaJrQdd
XNAtQKnTtXpmeYPbeXc28bjDQAtJABF5f5Ko9vKY6zeV4+iS7w8EdDHd8xjAIl+oQttqidBFU59y
a2nnTRA/vd9ccxvLgh7PT8JKJbe1MAKqgmzmU9+uUgJ40nrhXdmo77KiUy3zpXv+y0Nd6FlVlUgN
s1dbaVSlOOG2F3p/Q1JSjAr2IASPbJZYEQK9pC4Gv91Nv3CleeQVf2R4kmK2G08YVkBP4DGkE2Ad
Qb1wYwAd4L+vnM9TsPYhfa6IB7i+ytwNAxrSN/3UOWLbBT1kCTnkDSj+7oRTPQz95Tlrj1/u3RdG
C7uXkUdA32tyNafLcXoEI3hwVbqzql9Tjk0m/sNzcv35zDdgL3U1AssCoeOBOnl2E2rkvaluFC/y
Bn9HkJFoPNcu8jmYa9o1NSzeQKRcuQryC8upDx9sO3LOQWr9qTaVoNKSNk35bV5Mnd7HyV8nE7/b
c4osIxgs72DcHDwo2Uy70J4wX4eoFDka36pBjdjsL3tMgpSpuDQoWou3CCQa9sXB3xTYcEWsL83/
/fQty8avBmNff41t7YlZbWG8WzHUib9bPCIyqCuC5Hhq7ejTx4ZlPHDWphH0LU/MYuvex15ftxDj
f+aY071t8Sl+VGph78xDw2bsnvMSoSVEzlHJAIOqMqUAQhKbp2hcATIDtqw4iXKe4VRAkfuld027
jYn0nYJDpMqo+Zu8uaTCtOpgywGucVKXEBj23WkHnB1cL07D8SqsQcwMOlS0eO4kgO9UQ5MtpG0q
2rXhdCNscA7OSgQxoNB1TbEjubP4i9dr5pbw9qcdtP2QxdJRRx0a3bie9FtZeHoTI53ErW8/LPEU
5ikqHLfOuUdcNTxEo7vNlOM/PEsll7sEWfFQXv+y9Teq+u9XZc7qIXnCU0gARGj8ESG9hp56k/13
z+1orpIlAkjcZNDe9rg+0wxjz3ezaRp951Mx3HLmKmwUEKgFmvLI9Jy77yk8ub3CtoewLoNNz1yA
NZbRswai7+I1y3tY9XGgB4Re+He0QA5ayHxNVMKSy4KbyXngBL3433HYRyIt+kR289iOli9Sno0x
XkLtm3NzDnCktfopSDESUFWhj2fNJREoXtU0sJLy6j6AWnLMHg8F+nXW3vFoKLv8/8s9qhy3NBp4
QBW0eVqXoceefaZ8kDtmIjclPmQo0vtGiYGlH1WFTWC2ZYLBm4xqNrCbgP0tIQpv92wl/JpnU25E
ugBtQd2ck939UOXMhvWolSuZvTy2jKaOel4pK96QloO7e5M7uV1rufI2ijioPhC00eHmudLgYtMI
+Lzikwl+r+UYaAl5gTqECriSByrJgKosUmxAWM6Q9OAe6oozE8qy+yzurTy48LnTOtXEF5esaCv/
hYDcDSW2AFm5WgyooEPd7zfybTLfedlXnbnuuuYy2pZGwY9oZDC401QNbyvyE1m2F0CY/VFmBfqy
qxKE+jsr504KNPtvTJTHbGOpuDQqllm1MaeSKpuTOMaIn9TGuoiu5tt26xudvWVusqkdrnQkbhuM
6XXzskwUt9FMvxiip29YYh9xZb1pYpZjctGK88AWwU0t8bAHqvHWyeRha+DibymB4g1HWUA9AuH1
mQCgG+/TOTTVfvOOUKvd33DS8RXidJFpr8It/7ohrDxFtgC6Q06sICXcWq2tSjxF/iv1jRIlxQCb
fmo7CCk8R8KfMeoemDcE92sB+UUUBScYZPXEn7Dd7xYulSC5MOz59NTk1IHdg3LwsGKVjZ1jJbOY
RekBWmLP3owqhvfpMvOfiQQrgY9+gofj+21fTVYBSamJ6Lb6kY6mmQc0Eh1iB+Y1cugnV1NhfJMP
ilmM+eF1maT+yNbIVlVnJIsVfQMs5aZTur8WeY9yLTU/P5bYHreNehlJiu/+z9vyU3f9PHbtHnYr
sZpaM9qjbbXoLgQlbQhQv1F0sGS7JCuiqu7KqxsfhuXljuSwTWLlqskT6ceYgLj4oPtcctiBBoXj
YXgcQHb2BM76tzKMGQrwbAOKJVVHQjM36RgLLgqjQZ43lglWqF5HaiZuB2nhlYqpC5ezbpYtC8tz
Ty3j0Vb2ikCrtlKPDn2Iw0HRKbvxQX7+DiiguMFM0Hr8WITpiPS6k+0ogel59pXnOLzVEt7scciZ
pc97F9oQKeKNva8QVT6NvSut1EHV0YghvTEIiicYT19+scOvNxl7Zwdx+yadhYAnhxBQcaeG7dzA
msxhBaVPTFdz7+0AW/swYc8eZoWZ/H7OGo44F1q/gQqGwjcr4jJEoAns5OAuSQ8YI/Q6vLpZnB2k
o6oPZRuPmOStXENJ6ieFcYRacKtABXD0F5e/fXd8bs9frAZVTsSHlg5o7FkphzGVNM1EvKoKSAfc
qqfCjE6WymddFvn3L03FdXPilkAqu9pyLjAU7n8jKvZn67+fy+PaoevGHDijsHSEdGqD0ad2XXUU
9CPAWp6OCBmsWbpir04z9BxHJSTkKBCACMGOFh4TeFZTJ/qn8IAJVGGnJ7cSjLdJhQ74+pt9lf8Q
r+4V/K0iasY/zvqWra8hnbzKeNygXPTyahP6wD4mHqENSmm43O7TMx3OS0AhJTRTdtMb9Ckf+Rv7
ae1zXwOKpMmM163RqG0xtykYCkml6UwhpeK14C5HDJZUoAALWEzvp/GSg8x8JVdV3LTHaa8fYDKx
MhcnkA2PBafWroQtehMtYGZijXa8KT5/X1v64YtlnQypggm7AX0+A78xn5kmzalkdnD2Gb48beK/
Mo4Fw48plKt43u5mo1x39sNqzAJ1bdwUzLqXKgtDhzHV2z8Vp8+DHLfsrnfJiNPkTz+HhSqvsJ9x
jYlqOfuCt8xwyW6lpFmo7vBVp2M/Rgc8WuAu4kwfo8/nrY78otWktoIhHrFAHkyKtUA2ub5IeOXM
DihaNuyCLCSZUKeNu6wvpACgxzkQs03NVZRFJg726C9Z3v7yJbfJotT+aBUxwfzbyxeKHKRUDiWF
cVEF8eZDL6rLsroh1xn3qatOaQ84vgHpdpz+Z2K9ENiXqStvkxX+VKM9ho1gPzwhpuJ5SYlGiBV/
PLgowJygyjqVo9L1vawbVvHN2M2/2Zbx+cYhOhn3nGH9DgTEwW0poGbvW5SasVipIXNUqyec1Zv1
AdECldhPqZRi3ZZ1sYClAaVeR668NliH5AqaHQ0zuCyKTyrPRRIfQXlmFrzKb/9SzI/8MGn0YzmP
til+uQcb23JyXxK4WHEdg/gHK/atJTub9wm81p2G9rejY09+ZZLdGAifukuOJx+x4iRyHGSG5l91
q7bpnYMC1tCimHVmc5OwuqpGlol6g1mHj8AEUhP8FbOz03eKixVso3uaAMo5ujZTEp980orNm+31
dxMsFVCXJZhyVh9uMZg+GSvNqrfcV4EWKA+W1se/Z5xP/8DOIrlpAhznMrGBDAA74zfPR1hYMk/p
p8tBg2/gsyPlFRb0vUzfNfZt7mN6Sd/acaleOfDdxWofpp2SfDIiPOBiLGciACjtpqqIxuOSyjI1
wEeydCwdgMv00DTg+Ynuf7PPV3KGLabH4u9h+Ws34Omq6H5cEGAZ+Pkp+cAaWW6486qG/OuOW2wd
o6GuCtu9n0mcw9rvhJjUCyfqH9CHzWGEDjpQFcTJT2ZlJC/ct2QBUT2us/0/SgfnKoRgw7s9vLxO
uvu08q9rx4Q6AaDxLB6mDXMNDvWpRl1fxcCz6aOGNw5kntxnLXHLy1cjYN6VRf5JO3LNIudCMzhs
WTQzjUAJlVC57Vw+LrvOkrHJJorhnAbHU0L6hTc0wyzNN/yUPUUbB0mHceqm/EzoCKsV7P00G+54
fFlGQENINjg0mWo0wq7TF+cAi+un4WqjOYq8WHw69qFHvIGvOWlZM1CrEIHTkaNBY0ZfnudBV6UM
1aOfeKqM7JRNgRMWJ8CKmQwCNxyAa3YJnQQpdBUVLdivnQlCevXW/HsvGPnvTySyGpqvYdk6Mry7
hUfLPwOGPatolsXyYsSI4zhc3HnnachcILIqm3ocEO+Y2+3d9yBjIaqINxok4JrNKvK9EotbqXPs
26Ya7TZfcGCSrDG+0++8b24j0Hmi0W9fxFv8G1IqO3KL63jV8gO8T7XxyTGWPgDoTgkOtzjf456a
M4f8E27SGmTa/FegQFEzYcsDHlwISziTpCbTNac1jObj3XAuhaYNF1skkLMP4/jS9x+hWVcwxPsq
A2ZOIcZehCwSwt8acvySBOqOmBjrbU+u3JMEg5HYs/f+TWa3p+VMBq22UMGhjhNqL8fsH/kpTcvX
Rl65JOkSOqskXe4rL/6mMrWKwCDjR+q8KW1qnxhYcP121M1jQrBHdb37PaJLDjCrEKA1udrEiQ3p
ayWTYNz9TGggDrmMAJ68NqSGbilLykjuh0hrgD9rW9be3sKcwfPE/cIYMUB255/nRzJegF+4m8Vm
JJlaye0tytYG6lazsoeyL1AJXIhFPHYe/J8GT/o0eHHD7Nj12QNt8sLuoO4NipK/NJ5qIVw6tXk1
zmlosuhjT9pf0C1pkliNMyuqX+vBqn7Y5Wjh843LC4MQSxRv49/cHT9NMbTpY4KZyi5kNoUUg1Cm
+1c0W4PbVmOSgA4M5Ft0CQlxueDRbr/YRoaTG0IyWxXzk0DAW1zbgsHeo5qhnt0j4UYsrj0bwcdX
gGV4xnhYOS+6+8prUqvsvoyOPTa0k6WuZO3x9reFG082neLngYf4BuHS91hayfWJk18Zytqtvr18
edDaHZ15nlKkWP8Q3AosiPyycu4VeBs6p3y7gDHQ3yX0dH6uVlivsUFYhs3TRHHCFMDXuNYATKdv
fbufE9RhtUSO21sIFXz4XaWUeCldff4c5uX+VAcjsYGZSFQrp8Tlyg5vjhKyqmt39ajcJ/5Q/YB3
ut1f0RJS8hDGAfmNRcAmWqxOcSrctxksoY/VBlGoiKJ9tmjsd7+tA6iCjFshLkmL5DBToA36oAhh
Jz3WAdFk4gWE2c8DAH6R2/6Ii9R7PTAjFc2YGEqzFJmxYtYDWB2KQUgBi24kg0MFE0TIW1WfihwH
8/bCUwT8rWN3+jkGhZdZwO6rnAfTKx5kMJLGNGmWDALS0w1GDRquKEl7ObWozLEnhHCAG4yZtUvr
zg4AsleCplq/qkmEaDpDyP0lAKE8jRWLi4h3OLr8ZhgQks8NtLhhnAZSFfWUZWa5foCdE3iA6W3e
muipa1xHDIwSedtWhmDcGlUIunnIkteHmMi//TbAo8kvAvqwjKvi2JVwZgnzTQK9qEu08Mm55PLQ
epIQIDYfvwtBhZCxHgVEeNoW4cNDStP07g/+rn4fpyv8MuCjy/l1Nx7olF30MApOj/5mSEKy6K2l
uxVk6rg2t4ikmOfD2einmcitKbuYWeW6/M6FqzTKs6knZ7m3fBmVzc/0qXVHH+Diz77plcXwt/Y3
sil0NGN7RrpMEyNLGXLk06ej5c1gmeCQU6yfG17/J1ejo/4X5OEVPO3a4jQBiKw3X5yOaenUzr6U
khtREyepJGdB+Bak8eKMUg+G1inyOAu48ZcGtq+MqEiMtJVZHk/GKCmtMM9YxYWIE5pvJ7x4L9JR
L2Y77udKerF9Ux235XQXx32FFMQVlFKOwN2L0CB4lPGyATQUGDvz4Wej4rH2PKEaDvUWzbgoW209
KURoK3ITSr4Wb+RCFGJi/FRNsCRoI2vGXPYM5cHoCakeWVUCJWoNP2wm8yfcg6ThlYmWlQywVKIN
jWZLqh0dcJmJ7n85BzmP8Q73jZn9MGmTKprwDxMEAW1TslHLNAB3H7sa7ubkcsNM2JvBrtKiEdsS
0SKc0FurPsdBoPXJ6BXAt0CiiMyEUUDqEj5Pff9Rqdv79ldy/7zKHYtQb5NHPSFZb4Q7kzzQ6Xej
IhmNpBgMB1cBzbPhlEs6UQoualId5zLEPEz792PakNCzC4MMCB5ymUhY32fKVe/ybzI/P6BLyoYp
bOzdyjcN2sRGBkyUcKBxMSPYImggqQCIbU05uvAUHoHRJY2ctIP6G5/8Ytmoc90d9ljIGualrJAG
726MTxKorCQeyR/fODpayy7ISW2APG+ydBoRIhSbNlQha7KlLBygc9DCXqHF05pxikpxE0qVRE9x
xdPTntAywQjpNuBW03jxLbkGu25423k9r5o6aPd62q6LsMfelwkVy4Nb8zg0Heo2rAeTGR6a1DTG
npfAo7YQxyo4iGCGDvac/pW5PNszT4/oPHy6w4ELcF6PkM0PdbTqQgNFuRqESnSPrkkhm6uYt4bY
b43L5X7YLQ4EYjwSOvoJjHtmyk/AoWzEhpgC+UbWjZ51eeRA8ksLsdBxoYYZ8mqu5M6ZoYmTKAht
KhSANaoPGfx5639B9U9YBnT4BY9Up0dylkwf52cYoIPBbvELA7uFVt43utBkct+OF6BwaAA0dw1B
mndDRIl7HpFILlLgCGNiBlJPkbdcRoozzxUQOApp/CNYKytLoxZHlxmci5lAvWduKDFn0noqH8NX
6+uuTlIUP0eDJ1liNa+FdyOwYBTZxXsEDSZWX2On2TKl+Bf5cHFJSGFqdVXqsNxpxUuwJw7Dc7fR
ERLGbqnjSNAZNz6/zjt0qgDdCcTPkgny/z6sv6uBQWBPnCuY3zAS39NvjEErOCOKKjMOTTsY0ug9
dK90OFb1OM3qtybF+ZS5Rg3SKCRIb4V57eDA9jOBA55jQAb6lig7jlzkEOaJu6QSOHfiif67Kr+I
3eexU+paBbhN+5QArYL8lMCyRtWCEkWMIoCWCQN4wpz7/pXJO6rE/jW2WJQa2U85QW5C93HZr2e3
G4IwAFTN5hjNXkBfAMebUBMpOjzDlQFIeX1xDjX45y9abH/zeIciRv94RkSpP+vSYHu7sFJuAAGT
+8VCKCrMEuUjnIdRYCasTx/vM5IDxfyQKrXrK4rl3IV0+jCgH1QWd8w+nJgXFB4LHxSiQlvpUU9i
OZoaqCDZXEdQs5Sf6E2/SNmTUQLEXAONL46hskdLXYQnunjxRRo0dpphEDyNK6lA0Z5ahexVZaHo
bTk8ydFKg5Slx0l44zuKEt76GydWDRULrDe7Onfb/s/s13f/wK7V9W6H3hwLkqYeXqKE+q2Z8Ias
z1zwZRci6nX/79cGI3RZPYYjbLBiDSgsRgBLSDqdyKWQWEVKbmPBn7UmthskWAm3mDGT0Eo+oQrT
jbaSLFBIMTmAI7TGorWxAutKTIIVu4BXFw2COSSKkKA0avKez2iudacNdgity5ZdYtPd8zAuxsnQ
xM5nFJ//FETphP3HUo+YE4ExMI5nLPbFH7zKqaY5KtbDmzAD1tB/VLz4BzH41gN5Ek9WgoFogkyk
QqTCydaObbchY5KoWz9KSKvCd0PjnNi/V4NyN92BMiSw7KU85Rsb6DvCztIBVUE9YnCo2/FVL8kr
Sb+fsLZSww/wDU6DLG7+VJTI7VudExgr8IdKhhmIO8vHpsGBWwg8cYT282wcNdKdbLFlcPz65svU
xmCJFhz7LGob0B+o4gxxsSNC24Wg7pMs+dFHxJ6eFG/ZUO6ufpVEYuROUryBG9s/JWthT3ByTSAM
gCVFYxOnDev2Fryw4BlhNH5GF+u7KLTR4Qg4vJvHFL7L85O5W2YP8jO6PgrKWFH4E8j+JSUIZdpi
9lz/tXXDmTuGrtIpJReZ8b7xZrnM9gTK8jGb1Nvwb/f1/e6N07G3EgYeU0BWpGnybmxzrXW1W4h0
K70hpd1Z6clBsXiO5rhZR4x8SPBKTGfSbvSL0vZYCSNUDeUybwaB0q3EvmALbiptkXRGZcvBFXJb
Zn2c5SmLFw1CJqBXyPxSL+c9uWBz5Sm7u68dxJVLbxe8QKnWRvs66FIxJ1P5oYDV08cWRxH3cRkW
lsIg9UuZRpG1an/RJTWyi8e5TOE9VfiDjYj9/Bl/sJzmfX68o4bAwP9SYll4KmGv13Fd0ovQf3mY
grZlJMngp3Pheh8jxZniLrvn6KdpeFh2SwivScVLCFCRcJvy3iZ5KWIPOcsjsxVyttptlZ5vlde7
h4vfAcCNzlF6WGgE4e728aStqF7VWX2Q+ndr5PjF65QrpSkkWZuj9hqBEZKU7Iq2CsGVundAcyT/
qeaiUmPar3Jj1MVblYuqXiUbbXtLBbpURbQTQeZxRDVlUuwdmSK/hDT2uVzcgXEK/wMII2veBk4d
O6OLfBxNMOxDCjrbZve2o8tArShXXgz5k4MEK37cmYI6NcjEYkwg1Zt2MTb8X3mUTPsCxG9NvyvU
IcOT3yyyjPjh6oyd+EdL0hPQticZHNfrsMwZM99dEiVgO8Ub4r6VCOYU0AvwytAXBXqehF2s2dUc
cLVtRVuYJz84WknLc7p2TbMgSNsBlpxZjDaY+Hop0fxOxk7LRZPL+elrmESISk1X67h0ztuna0mb
NV8v64jpEzRHWM4xTkWCfUebLieiMqZScUKkWnDUTHHV0SnvItZY047UZeFoA+T3kx6St0yz3zrR
uN1xHvcnZlh0jJ2Cm8zGNYJXXl9ClC5BKcPD18gAjh38/1JyRuxqN4AX49qHe7XLIxns/tw1OdWc
pQb0z4VdBhdCs9pLzSbMcWREu6u3ArqRQ5ly04bU2Yi1cf32KohmTapBpQeXJi+RyKlpKJXgwFVD
qD8C8ZAXLxV7oT6EN1Crcq/w4GSYG7ffHGa0kgpMQhXY3+na71yXK5jNfLm3wWmbbabE7OM6Jqw4
oDtc7o/b0H7tcqVWy5jijPPIXZklIcLGo70SVuDbWqckVOWl3RZGMBr5mFWP7aNigJzRRtAjN+d+
EDRFXzg+Azpu2Qr8HksIQ6M9b0naHR36wD6PPtsSk/p4NvkLX5q1+NbYv/xMhHSLwI9pjlAtmsU+
OWsDxBC8LKFSDAXkbq2mUHZLFDrfPtUFkJQqlCXu39jdX8wPkyw48Cd4CxqCrN/0eJVVDhW4Qrwn
FAqaoJJBeczvi1luCjQ9pa6AKJY5T9Kur8FLjdt2m6c0sldaesek7qgPNjSajDTtuQ7G+2atSYpl
gCC7aBjAoAnNLaPGyTRYmIdMC8MZXXikum7bBxEO9EO5Nphnk80Gtxbydb9fDQCXItsEZtOsSq8n
r6klZrBOrSsBOJPq0wiDLK9Vxv7rKXGHj3W3lbok9uJDS1lavOlRzY/o1LV0vpUDmlZpCTScGL83
dwVJVqQ+MfkXaeAzAWomayiajWB2A53Avf1f4WBC3Y2fIGuqYx7wsnUBTW2RusOOrsWcac+XOhti
zJeSI2RsHBeFLe3dIJd8oPHgDS26DxmESnr1e4DofyzsrNoEw3MlNqIfYW52jLu0dd3xOlNmdBhE
t8XHHRD5aRNDabKtbJgRLsgP73cJ0fwoAzai3L6rlg1Pq6ehpEpgDEflmSk5d7+nqstkND1cH5qs
5a2+06N5zWGL9GAI8IPNiM6lUcjA+wmzx0HDns5uRtFtwJInuivCUv3EuR74rWq7Yr+RlC7LGdfN
zkCcdXX1thcJA5p2sdT1YLJ6wJbfRERHWuTbwa6wq83D7izWImxXWjRln0kb8ZAtjgr89TChTQbl
sHlMUzXrY/QSOci7MD+S7s66t4T5jG1cJnvtpBNnfVa9Amixt6awcPl0LdcYbNgvYqmYjEyUeQLs
QVHkVoricLmm/wCuzamY0XVRLoQjbUGCYKYEusygJEaLYaHjGBzrZtGBcSNuJfOTXfarJz3HiVDy
ocrVoKlb7KC/swoVA8NtwFe+AgEfoapmO+Q57vbkPBO+0/W2DsJU6hS4UaxSR3bCFnNgIxYK1er0
Iey0p6Sa047FRKRCvC50tTkd1RUAy1lR9RpdNZad7nJz6fKM+xbdrdjhyjwpLYffSUlBHOSobLI9
qsNPpny6I4jCslypEqXIEWyFuwnIoVfKBsEt2XrvEiFqF5+vSxVbb7J0pxNW7ZOTRbAqOxhUcb0q
/kNP0k7UBWAn/JJfRCya+nQFKpL3LNOUSZ0qw4haGEWdKYkA7npMox0f5GP8iovx3rfHkAsfvqSi
0lKuOwb23v3I6WbsAM4D2l873EePiWF6hZoDtwf65E8ce0XVQ5eB7TLpaG6jBWflb7yLEML2x26c
ITslWYq5HqHav7LjRhroONcJ7ESx+nBU5A8/v8YfWKu3vHxAOWzgFwJAhJ1MeQIjcULkePlXlifk
x47sjMdqAst0YfRSyj4ENHX1JYUhtU6maAqpmSLXd9e9/7mWr48uh9uN8JR58eiWwNIadpd/kuz+
sLQh3MlldeDYC4s7Xq1cuv6WSsi9uDHX8YNOX526koYleHg1whM+rHt/kw6AgX86IQ9wsyMm/QIV
HGI5ioDJyn5Ql9FiRaR+e1JRmAy9lVUBNZK8/XNQjReZcvqNDnmjuCt4h5cYRol3t+yRfJofoqOW
5QiWbikPeTRN2rHZaIwe3Hj9RJJtiHvBTjqfBLmGAouvk2fDveA9tPPj3Q3nFueK2KPtaranBQyi
6DJ9I+975CJ80upZW6JuSBGnYODSHh84miSgKfCS7fagR+ULhemxXIwMCPgaIEevu7IH5CB4Cec8
8qwt+8x+26sHd0A9tgudLLNIzfC/ME9eON2p71vr6I2jDcC+po52XtuGLxg5XGOi8bNSX3AxPpRk
1ZcyBJk4K5oNjdZ30QgqgukKpFnFzl4PvTLJdCjyEYSRZzXtYUEVnp+1SU8TN8zEkHx0VsrdxjxN
9OY2NUyCqI1fdGINqW9K9mEKFqF4fyv4kkgiPc4XUmI4fVrt9XV6EtoqYpMu+FHQlP9yQa6PpCDp
20Yhq8uhY8KhwepxbrhzbmOwXF90jHE7245AK27zzSo8P7hyPZr+mFF5B7vhZCqlvN/+0FfuEGgh
/Q7R/gV7puPCR2BwszgNCClf3TC6AU3Pegt+fiY9Ip+7qGslSw+G2pjX6zA/TIy9cdeeYyotjgjd
8nLVCcMOe12VEktmrlUffkAOV5tlwQUuKAOhM+HHL3+hKFcicUmht90IA0vZQ2CYGQhJI6N50fL/
jTqgk8OcOGMOsbcCJS2mH/ovBqd7KfBUbcGAjlsE0LqTQoLga//S9QfCcSPbwE7781WTbd5mQWhR
yv5j4RABj3cUuScCh3CXU0pjH8D58LV6ZiOhZRX7tDK2CgWOx5zhwgsy6Dp7Iy++uv3GGOzhgbu0
gXZUKD+kdBanWkaBfj43NPj8rdhR+Rx6djtfoypkVV3vHq39vTwN3lMR1ckdY7pCSMk256unR80C
UTiTgkXa22lp4+awtVS1Wp5jNjAnxEFwSEW7YBmVNRKJKJWu0Kjvg4pGz0fWxyfqLRZ7mT+Bj5HL
7AOGpqPx0GqycTOIK9OLULh1hpf3OaL/JhVYIR9ncXN7+DS1LP9qYZ1RfaC9QS/6YmtABB6WTADZ
nThkDjNlcBsOfM1azqXYs8ZhGW/SxyB4VQk+H3NUZjuuyPkg5nmwWfpLErg2eupQzBweBJAKcJI3
B3nHwIvJ0nu5tL+EFW3+49v4Sky/Bl180olUG3gcJxr5umH9aU2i9gDEMPhgEl/xe9CTqjPoQ6jH
Ga6/ndMt2cmv1G0wm9QXxJEKec9mcHlDeTZjCYfGzkMsfLQGFq1VHkhwF3CkVit7yvGT+JXaaGq7
kp44ynhBkCOI5ctjyKVtQ/97xj1QqDse+8mnsKhwTXYv7TCKt/EtN4bNUS/1mWauNz8kr+duqzQo
ioVK+wP6zRLEeynjiVufBDoNcEpanzE6jBmPwS+XeteywTuywK2TT6BUo+wprU3qUlPtvNHf9eR1
s5WZ/ibQKHBLn2PALcncXqqYVf8jA3xXy1LVEWwB6BSPXSg22fTOtWkWKQAEd90KlqEV8ThNI3JZ
JerBJ12Czd0fvlTmh/qDJKjJWSsdIzjYklKIv0LE2vZNK/zkC+AXZVFOCI8qUi7/iKf+MFiKHzJe
9HdM3c6HL5ym9DI1aWAo2XxEawJR3XOtEeRMoYNwXHYyaAI5SbxyWdSjKfrMuODEUTtEg59vyFgs
AbwlonkP41vJC8D07CLEr8WIM6pKyioQrqxe75yqN+HjgcYukOppQwPhXV8tnsVZQ67cJlIgVYDe
gzqVQ7jURJfWUrYqp1CS5x+GYSezf8uhoRCjE6VHfdbZ4NSnlkNQbtiArTqwqbqB0mMXdI/Np3ff
SlOQtOwE8MhiksVNBEsHXUjZDZtivSzfYxyJM55dVeEz6QE6YhJwLTji0x0uQYPnObtRGEByDcKl
Q1f8BRJ+qTo/JR6b4gv0EPr/89fF82LTmnG9F1/v/JiN/pDBt/AuPDkqRDD6XThWL1HQB0Rw4lLU
uGo0wwApNJTkWffgpzwgADv2qfdum9OH/IDC8+6l0SXlJs/NyboHIBPvkXDacG+gskfYQXSfZOtR
RIu3u5PEO7qcvCtbT1R5CN73TYlgrqAL2rJIJ+mQ8jVI2WsMUrBVQEw0roR2LabhpBfTqWZ8hRl7
k5nF6gaEFVI2gw/0xZmO9PbE7wcX++wrJhnXZ2qY3Z8bRXGrdwv2ajM9nkbo3CIju1bfb23amQJm
9dcRLS7U4aLFEtv/UVXHeHAoWM9iyORtvw18bFEhzKZOmoIwSwT7vv9B59dzficRhjjJ3OlJbahw
RHkDes6mGr+0L1s7kO3toLm2b/E3GN6AfZg/WPJiUoXmw7PeMN2qUtmn19sg26G1nyMA7RQB2A7/
25E0OVLuvpe+BNVaU32hmhVHQK+8bLi/h8VZALFz50h2HSCPyFx3+4l7nUz4Xg9iT5jCYVVMdxLK
cKfe5f7J5zYX4d2MaTpdgfEYhHxcfsFXtuLXkEHbGpysieXD2rWjOBRXWHgeq5sRYEPlENU3ImUC
LNGdUWuAYkzrHtyxswyO/WAjBlNDX3haQhoxi0ntOyOp2UGndYeSqILrPqb2eljfIUqbFY2SHxFA
fhibOP0RdlXCxQ6W3GZyMP5XbUuiL/pTqqfICivoDRM1ATf1lrCzFeTivNIMW/lq2eaNErZ0RgMz
pP67RE8Wibr7i0XZ8XEexinDHWYqh6dgE4iuEFZOSk1lKCetDpvAkY5fAu/QewdE5Y+U1ueabMhy
io4v/3xYWxZyfKUaEzvFj434zGGR0TIYPQXR5PYoCsH+XFe/3Z8ndO4iLWNmOod3OXyl715DjPBj
T2qF2gVj7DQK9r8+/zkRkmY/zbN7datGO+sub9ZtYZrNdDi85vWxOrDWLY6rJHK349p4H+wtekLJ
sg2fxHGsMTlv42+qtFNKQvoRHIqHx7klNUVJn5DqeQNL7zvWPSZvbwsHkhOfYQQ5CK4KX0k9SC7Z
upAAqz0yKFJRwTIpv6SxGni1SAR6sqWcaEXG2E23HKHeZbIekz9mffoDxCaoMpNLoCpEi2fvlwtK
PN22v28d8Dgxv0ejErzhMr+vE07D3qd+c9rfNnAM5KYipKdWZeCJWB74JYWdNveIG2yIoGRpE9Ke
h6bliaRx5t464YZUVnwpWOJUASgf6JLWnOVThUza3yJPX2pnggSEupgqKYb4YimjVnwtyRbrY4m+
+aDCLuCxN1ouGhacVbT4t3WDiPgQlayYF9DXyqAia4N121pGw+eGaWt9yfM9W69mcyjZYHQdCZP6
FsgmO+ajBPfZNEB8V450lbl308CWB6BsWmIJ+SajGpj0wgkTKk3/Vwtuf/PgnTx+EX+gHUcQez5W
cUeO4Fo+8u8FYHW/iyGRsorzpL6GNWrz8zmHHhQJj0z1ZK4PyEKtprit1CG7JfnAjaDIdDUyqP7J
sdpden7/N+6ZLWXZ9xw3nMIaPRpUYNNpEJwF52Zl8PxXjAjuszGpZQowZ2AH/SsAXXQgsYZu7ABz
hteCxS23PxKg1p8zQdpJcj27JA94akREPgDQBgiV/iLpGVKxfRT5u6f7R3uRp6HsHjI+abWPzNTR
CbGD0GKKihrGqG1Vx2ryRD1XrfWwHQ8b+/v2uPBZqH7Q7Zr8x3O+w3fXBWrgZHt/np+KIhPJ8py2
vbmNYDLWgkeZ5fU/42nH6uMm7vU9dujcYJpyKEQKcZPt5s4hGJM6Rl/xw4laiQ3SKfLgO3XFNADh
Wyz6JAYXG0NGp/1KVdQZ6pGBT51ODne1WTouO2eYvd9HO80oGejUGIxSsEMJj8Coom7MDzrONaki
NKFlYaZ8TTkLAyG4jb05KMZxOulNYKTfEJX16ihXivwxBtF7zMbjSaFiv6IPDxxOa1Xyse8Cig2Q
H0CEfx/zdvO/8H9C2BHOvDdswMon0a7k28To2yvnyzx03urRVpfzYURpXDbNC2vINxG7uUNxSRTE
M1aHOz5CLQ91PWq1tS6h9gnl3Jjg1Kulm1i1WvvdpukW7zd7DT9E6npIa+9c0eSCPEyHoNYaRUwq
8enSn9Fs7wELViC2ryCo3mEXvAmICEA5IHrzUXp4LzT9XhJYylXNwfzBcMRjXkpAVWocicG5LCtY
QDIXxCGA6ynU1uwytkIdBN19DSVxl8P+YpwoQflN/nr91uVoD0PHXabJnuGIa5F0RmN7oRs1rB8g
ZMfwW9/e744ACW9R5NRfcCrTg15lxWLCrz8cxPXEmrJVTZ2995rvXV4QKKf04CDeeki+OJ+g7B4R
BKgS7EIoJpmKPrijts4QsSi0vkULqSRWdh89JyIURUnFkOSPoDK6I42AvfYB9qatRfjBF3HYUV/B
ihX9V1mRFh5rHujMmLRmjxhM5oCutj7K2xWzcRngTavvSUMbdOxo8oWKUeBztvZGWUbkgbxV9k2I
gBMDs0cj3PFcdpVOhlL8mhS4/LaHzuJH8CQVuX4xBfMtCU7Ubqgfh5b3NGXGBdLdjkY5j8lXXkjS
o4yXVo9iu9fUFwM5I2CWUwuApsfzmIHyOvBHzKEs+SbqdGXa8sgkPCCsjrfg1oSfBQs/aTCwMqb1
XRsBaUtu4yzGUmAJtrkbBo6oNhnc3a0y8o3AM/7g9H9oYQ/cngzsWsPyDKDGvn/GiAftp19dU9Uy
VZ7Jhrx0mOklHEpNC3iWpjix5NcJsfFgMozqZKDNZ1QzIOgsRuktJA7PYLcvNpXvwdkpyZVAeT+z
SPiKLQZxZL8nxRnsG6JpKV5rtMzN5yXV3zk7nBKp9Z1OuWFSTTJCqal8B51uoGAisEwNnVBcDbTI
JY0nFIjkvefjMSu5YXyemunjwxGgxCRC9qMLIPLIgoSyx9nE6i+7/CquNnUq+gub91/cB4P9z0vf
1yjvLXjcH7xsdpmzysi7xJZJfvH9FtB0pZ/fMXA2kIxgi/2cnoioCruXzQWTmfXatO4YI/A6W2No
/CzxTKNALfWb6yT3DzWXmyqy9CWzYtn0MtPa9kbzWCbKjXdLMkBBFELWc9svsKKYUKelOvu09gCv
pbmvj522rdksJMBa1N06iwtjI1/aMufZz5SX+Ry1wworUDppKtuukqVj0anUuXCOlsNTJHA3ZBUE
PIT94Iw9UW5UfqOHJvxKs0YInnPs8tf07CIvD4eezi5+GEpNBiR8oyWsXVa75/SNrzLSsju0qP66
KWg6Wwcn0klIXawUw1/GVTD6BZA38RwGq7PD4s4OxaQXNDhubvVzuCMmgDvEIYEZ5rRHQ4+NypNE
/UkG+psLbJPAwHyA7Qb6SITShP+8yiV3iL6ZRAiqBbxYPAFmSvF1RDTrpOlpPiHipv1ZeeBoH1Uk
A/Y5wpTDlyMdU5wMZDgsKCstBtutq7QhZYsL9iROnAUatxd8jG9RLiwbiYrqq7DRH2fCXbQk6KzN
obzz9cMHxU71AnlALZIzVEQPgJb4z4VP/vc3kkE8SfRxK1sgp5J0hL38E9URtloB9+5ZgpQ9SUDW
xM5JJ9RGlOmy3N3QhckLHTae9tiUhhevVFfhxS46nRCy8891ggMHyuGlIgkEoBxMRNVdknuQdzuS
QYeStEevG65/7AdTPq7MgDgJrlkscNLi9bB6BhrWwk5fbgHxb2dm23E3kHHA4abMHgwo2R+8GZOS
86JOlHPbIxGgwOlJKDVO6N7F61keXx6ZL2Pq6kqfhUuxKjrUTv0wLGLTRkpeKSVy1Y8JD5I4Oix2
bfJbKOlH3aAM9si+oejqVlJ+J3ztmOkAp+WzyYbjCWCQCXuNx9pS/60c03B5JShnEItXf8lCIrD8
yHnOF9DpxiJ1dOdqDG4hpDnwDsK/dOYeR4hzjIUnxNBeLEk5pMxjm7Tbm/Ijn/dSVUjxsh/BMMDg
PDPJ9KWYdl0+px0y0k4MfHCmSRLQdtks5azh2PYaTuILazNYeJKNfdOC2s5JHakJTM45RKg759ep
4ZqHlVcWAyK0SL3pt3Bhj6hF61qgg3tEByhkMPun6Eb+T6yPuG+qaf3rlrH43wlTa3aPvpdCuvfJ
75DsX5Do66AsfEyOKa4oaSKKOcFldRZ63n87ges+Dd3zKNWZpVeaPz2Fyr+YMFQbKw8pNlj4Z1dv
FMbg5wLhnvyPU1Knvy7kgUAgeFCBTJZiPZltb/HTBbUe/iQVJ+oVdYf2XNukypMngIi7LanaHMpa
3xUY2Nxc5zrCqT/V9c3pL5lrcqCZPIVq8ZnH9WBD8m0MzhSRdpXnl2yxCh95zbGru0MyW3w8Inmr
so9sZqIuLN/N2dPvXwHoclKVUrPTcaS4eom2Io4nfLjG848mRmSl8B4T+0H5EJaFhSO2JiCQwqMc
FQ6/wMd7Et8u1hZ/ycSD5JoOLKCK9kFZ5/IMzvULTOLOeiFdTSN6h7Y813qY5ImVytkV/wEJbW5e
8fe9HS4ExjFEqrsGMhW6hEk63rMDhCWyN99TktEPdxnW3aqxjrXfrVOLIVGz93ko2Kf1lo1/5oTG
fP46g740IbDC+1diZ4UH5be5zZZ2TZHCYIImQ93ldLdmHZAXb3e++vcKptWaIsr8SASiMp2FnbOD
cqM7ULMojdNS74i4Wvaig+LWQm5yj4g0JLf1cgUFgbl38gGnAJx+f+APmtDb+poCbgb7gSsAvV3P
+NZO/ZYp1W1hmAZ9Wl4sjCb5dYptpvZApqTUvN2jZxz6kUgI7yDjOb8Em8A5vy7iMYJIz4xsvS4j
3zXuC/igC4RXq6fYeoAnGsnrEBzBNVQYJxY8qVXeQdidP1oTZk6uo4BpMeQJmR3tKI1mISZhSmIC
sHUV8WXrmg9lhHBoe3Tgg+++O7zhOkR5jkR8tBnu/E0Q/XkCLLRwo68rnLIwm1vP3M6Y6uV+Lklf
uW1GowjuTDl1Lyc5z+WBeq419La7ZmzYOUQUkwz3hsr3cagIPWePiDtCWTUsPSp03YcR3jgaT0nV
rqZUYhcIBN8pivszKh80uZp32R4lLAJ5Bn7rBtISMeRsjxXRLZ/ArseVwjNceKwdsp6zd4NpjuoA
hF0N968vnvl1RWBZSxad7houLi9FVSrQ+OvSdcIl7gfGEYjVKcJo7GMnZ6CLopZh3ZCoA/LWZ0bp
D5YM6hlu4daPumGb2m6KXThyxZ4V04TilmqNuPkgMBL8l2UAjaJhS0swo8qbzcwGg/Z/zm/RVdjf
6Omd2PE0U4lG8njiHDhDWsvkXh9pGF7Kp3kJ+098NFSRYi0Ofj3ZpZPcIQgn640tMbXSeKYoT1sa
y0azuL2kDrQr+jGP7E6s5GwixCnI5E08Mn1ZQrdc0sNCkajdRZ88aixXIzgRvPi7XhT7PeAI7Td4
G80weNDFGIZDvkoKEPv9aUxtRlaJy9L0MtXuXF2VzLz6MVk8+ZdkcXyufRXTEZhNi3c/uP0Y3sHB
TNRW7dxWGFgnnuxntd7MCy5pkizjYx03BK41EZdGEn1GfFVrd1rcjdyInEpYwijGWGK4sh3Jr3Iz
2ip3wNaqSQMFvxT68WI/QUt+bI2PVjpCb2zq9Z5CKSRdFbNohAQ/Ppjnunw+FtC5Xw4Ki6JhzIO3
bcIumWLUUGsb4lAlGSNe32ve+7vkyhITg1agqqa34i3V0XtI1BGmfu70+NoplzYa1RJq1kGoeT6q
KENnnqNp0rdbBVNwqz9ZA3vtwV3zTHNr1W6oqkWpQ3cPfeo922FgRXmf6G7pG8grblsUtmoqMTWM
FaN/1QhRVMCTT8JKhSQGPzekLasB2kCHrUgH15W6UmFW6tYQPr/hGuE8Pec5qOLOx73Tf6jm+qD2
+Zjt79A0y2TRLm+E1agRjLLuLxeRpX1rqI2/F2gPZRw5CnCCALKJtXZATsIjN+wgDBFynS0LaR2j
q66EmI/fK/iNBJTsmxqPUYN6rWVmCGTffnnZBIhf1XGK1OETAGgZ6jxPnC/5Fsa/7SL+ESZdpK2X
jQI80P5JrUd/p6dDyJIDDb/pYmCXi5mUOWhv6w2b0RltYI/L5Jg0JPyJeP6dAV+eAGT/Nzyhx1S8
LCAbB4YGtx6a/MDou3u07HDndTjv87GhMkOXkGvN9gvCMMVq/3xWIW5xyZF4igVfriSTwDzz25vf
1HotsfjknwrFLiejPLkAfnu5W/+vVZvSEfreR8Oa0YR1RJJWKc1ZfOikU5Y2iRKXFRughU5jwOdP
TtvpNaYb1f6f5fP2qYqDWPqDPWOIKCPPJzNtOsCZ8cptestZs8v5o6LiblLHE+N8bYAYYFicOvm9
kRugRXoGssxou2Sv65mcGSUOR5LjeBfh5ZWc9yC+UXK8XT7+n0bR21PalbzZX5vUSBxxVFZ5ODPM
wrgYBb8uh5fI56QUOmixMiCiwezUuWax/uP96mn29PrclB0Nn7SVxTm2k4AU9mghZsQS4bnN6wpf
ZPeJdAgX+kylc9Ujy8CFPA5zUvyUlQS4J957RmZijrxMo9fGeGe4nFxxwTiIPDqkcapQhuaQHIxA
dPgLKHLMfG/gvSmi6j49oYWZYuV7Hkqz0CI1C0+mu/86a1aRpHqwBTZF3aGote0t39/84iR8pM7o
kSMeg0VN+91e7KwQBoiBNc/NwhbuVmO/EdLZj3MSUZAQ5PHS8GItAIwwrTRmDHeW6lNdhbez0Kd3
sGoWKDjp7a9ahmg/I/u1U3CgefpRC+A4W6t4KsWAhSEdcIf6Z56sZIdGXkI+1mQIwUNhSyoRYrjF
PDKKwph3fYED7yYGfpQbKZQqaS1k+9pwHqqZ1j7A1fjyYx2WIFHtTS9rJfaMr7qmZmS4A4fw8KI2
DhxnMSWzB9Pw4HiYfI357FbRG3TqumZJee+Cx5k/7Box2JQk0L+8XOcoRywT4BJkBprL02m37sIF
yC2PyBYDa+C90fybupUU5bVLH4RN91yTYasx9qe8+7HOkOZbPY7jhduLl4eL7Xmh+62DhTpxHlTB
fXGZdvB5Av+lAZQ1gfJrUXm3W4KRzEaGcKGfI+2/KIClOB5U2IO5L/wDkXUuLX1qNIcCn7BR9k0x
9iCeHyYqzHglw1igD2QWGmxlNd3W3qGTbFvA+2Y71qKLeMplqb9TjbFFrVVhgkFMuIgjBtZHd6cQ
ISg2br/37HZ3CnKS+TuGQ3X1qAXfalbHnmUY52ik4AXKdl2FPwryDajbnlPglOtOEcxXwtamIf38
AmKxCF+eNz32iVei/Y2fr5ShSVq1rIxluZQzaXjC6SqVkjk3kJLMMGF6ORTKiU4zWyI6H8naeDu3
N0RDvR51jG9lrfh0ErdvVRwvbfBgRDjhK+zTM33w2NMHRe1dhbUotYINz+0G4UHtUIPGHwMULlY0
rxo8mPKTkd6FliK96EuJakp0tQKEuYe9VOLstDtlAMHCyUahdXo2FG2vhGEAIrb2zfwbwW8VIfmJ
KpR0ujPi/xtaS6Z+KffcUJE3DEtHC7Jgxb3TTHEgAomNBBxXX1IqECqDtPB8BfNVUOFHi4xx6mqD
xMSDRiKZ4gjVm3fWVQ0nNfQb+MnIdRqazAcQEmvqLdYJ+cFA9YSL7Yf+DpKcm4tmj1O0QWgWqGGv
/D8zMCJnTSFrEWpdimH1TJl8kazbgNvmdCsuH6/WuUX8SlmWF3H4B/Z2I05MHePKvc/uDUnmvfmQ
z1bgN33j04B0t1Fh/BUi45MRdws3+Oe5wElwOUmDa7g8tnlfEbmuTD8SzeC/cPFPxUcC83tuJ9QH
kC4PlGjyPR4OemwKf4xGMc3yOVfMbETVevp6z4cZFLso6LhlUwD6NbWx7Y30kQGmRzphowRp2bfA
PNurjTeqoq8NLBnLh+sJogw1zrgTrkvNoDTNHt8+OuFeCgdQH9tIzu4NhvteA/OixZ3EYqVTuwlS
lVeULtmccwFPPcefEvaMN3fV621Ef62ULTvWBsTFZm9Jc49CSGmNgxmpre+Cyl9FGS+hUBPhYByB
DvvO/NxXrwRTQ1Fg96I/J2HG/mpVxE8J74IP9bPNUkSst8RlKkK0FSLF276Rt99A6G/5/2O6fva6
+qw/wNI2v7chN7xAo8i3XsWKxpMZ5WFOhahMO81V1uMaTINxyYvrAOnJhGGMsSNIYqfR0DEEgq7X
a35321EkBtQ2d9URoyx5zKDJmWyyK5I6GEfehqWmPTkjOOEfguUDXN/7IZwuw7QM1pHYdZrn1UbI
2Qxn0SnE/x1uaLkMHDcRJBwOgYm4KgdbL8WYb+nCMFBVzRtRU+uGmFnDelmqdaw8uzCqnZLIDBwP
Wp/0hEhztT4flGbLIisuwWPz9xgtz1ZIEfMqg4Tyy9KXcCkrW3qOItVoy9uC88weGoTTyFP6QKe2
N49bPKEEpapPQ9iYsnCX883r5pcA2c9FPY0KSOV47qow4uJ3bTIWb7WulQSKmfGr/RWf9H3Ijkww
0zmBhWHIdtyXGWZGAnn89cmmsHmc9FDn7xXJ877hENzoAwaPV4pqqVJcytF3E6UaHII6AMbM6LD5
V45oYHp3IlDz7S1Tfz3kxI/u0XQWr8dENHrJcBrgPFqSl6MwrZRzKw4BV4CtDr64bWKOzu4SD8Cu
botVpaI8zIYUQN1QYsy0KmJeAnbSZZvhr4KS9/zVyUAZqcMJ6iW4E2cq7ct/vb/dqduAYQbV+qNm
Oqn8jDmKTgrSaT6qU0w3xJlnuj54d3E2AqxFANM6FH3MGdqFwBKv/JOY0BQE8XI6wkRIxzVfzupW
+vwOjrrGmlsileIaVIDQGjsCtG6M9CXgbG5O237ndSksgNW8sjf5rt4kLaU3x3mwB0q8ct6+hir1
YFbaLIbZNXLwX2SzGsRAsP852jeapZXBFY/07GuvWkyP/36p7apliQjag5tOcFtT9TMkLByb9siM
AksSZAa0kyDR8Ds8vi93IHQZOc9Hkgoll9pXgl2+NvVAoj/j/ec13r56LVy6xlkIyrSK1dJZ/OrI
uaNIe1hVGvp7VYhnSrCpEwjrCaO5mjkx7GgcO9yCK1F8gl99H6zyVpQEp/4+j+R0uu94kCug4SUu
l+O80ZWtkCrZjWwUKXviP4h9BZ61LoQoKB4eTqxajF3QQDt9ttxAtKiN1QRkNhUvUNcIW4IaWNhu
ZkCkJw9NK7U5IB8BGZUV4aRk81S2dFTxCOucKZiLJ++Mut2MxUk1HVaxWc5fSS0vla3RwHinX6U/
cp+zEDo1TIKe1Q9aLv5EEq08QHLnjHeWzX5U1ApFjZynO30/9r8xGfPbsczr83JD9ZDAav4pQcMT
Kob2eRmj2g8+yb6FdWTe3r8+1fyC9HmqMRkAY4W1gA9p0lWIrY5Y4dTX+KpCkUSMab3f4sLRYgKu
7UCKKhNLVY5K6U4mgTxOsxgqMiHxhUjZ5oI7+sBKJx3RNKwkW2invxBt7CZMHQmrU+9APdF9TtfV
ZU6aX3esvCSPbQHIcIEh30WPrzGh+PN2pArlVDnbDhowu8n8oVfHozkiSNmcK/S/zRM9J00f59BN
s6OSe9nBi3mMFjykzJvYmEwY2xriNq1nivx4bM6x1N0rgSN22bqZ+EE9PrAuT/6RgZUlghZ00exn
EYGVatKsHE63g8NHN6065vx0imSL0GFb1GKLAxpEl4y6BhM2DBCvyP3gxu9kryanhv6/ADjnYcv1
niISAkuq064QSZUSVRyqNnpUw3oF2oIWnDLlYhdHAiwfsgDuXVUQskt9EmmzAnOqUHH3Ima1X3C7
mRrDvfiqe+Kd23DtFEMd9xQueT2NwDZvOtpZjD9k86xkH5xekNkw+wfYco4YjdwWIERit08l+QCC
9wpC6kzdrYUjldXbM3zdve4vTMFlCiyrsIVHVWiEOwcvwb9UqN5FCFCgBAIfPEKFHCsrIrsPyM+P
gjbvEw0/ratoCWpiqgYqDWgt1yN2TR0e4ULbPsjtWNmCr9O7PaVbYshu3uuQEfk1UJsP9Y9gGfpw
2r/U0+gWsCB2S70u3T94FlElbHIRPV698JeXLRD3DA5Ii8/DXDNeOBiculLO3uW9BmYjQzUpiYw9
TT3JRW2ZUeZUn2VV+4H7lX6a/crKajJg3ZLKOPvj+M4PVHpnZNkZq3Y4jLpywR/n7RO9sCrTU7SZ
M4pzNzgpaIX9YVLDnCix2Uphe02FvK9GPTB6BhEzBjte/ymGAqbxjgPHUG/EPTsNhayFyo4/gZGL
yh9nEKmzNeS5UV9xusq8cjIAd6iZvjVB4YJ4Bdi75jCenxgOfnSGhnscWXL2arW/8bBlajSgTdYa
VtHbdhGvcbanF8lM4YzKMXtWFtBA5fhm2zgUB3b3stpZVrcjLxQ4XozPEpREpOrCDLa2BkPnROUN
NpqDCKRBSotduqsXnq6Qt2Zz1TimnwNpmE4JrgZtsZ24Ummh3xucrOADAcSRRqHQVj+t6jgPVKIw
aotlvfldnPtGIeVGdZr2VV0/0Kjbn/SkqWEYjpeozNOOAw5w97ED4WgJET7Q/goLASUUZaWD9SRG
p3pUUH28Cb3E5gvjyTbAuUMTS3k72tlB2GEy43Vc1ARzQZl5r28JEMrUQmk6DGFzhFbkHr4j0PBe
gU8A6TBOk1lcfgxjlZKxdH5s5/kH3Y9RtWMdtNZckvwCLVEX3hLLzASbD0z7697UFwyNcGCzNc8l
ysGuMWVeopoJZY8RmFMq5fJawmZqdtZgrXS1W11lYuLxZtMo6DVqSv2DI+qx2TPGQA3pPIP7dItG
5bsriznd7PWKnkCYNmTWbxIqlywJJlc2FgfexVx0Pl1cre6H9h6hGSLb5cQNRbSfPYDMhyX/Gegi
44BeKwufKjRV7aqpIHQ3AJHnpjI/e5ryUtijcpxw3ay7w23sQx6AbVRG5wnMY3TJnGdFD53aQHk1
I9j4cMahBNatNgWzeFyY0s+RnVK/R6gkzUynrc/NkXaIqMLARmoqjvRR90Ki+Q4TtAlkpZ9CBU0/
ahdiqT4WHIqSquUxCfi119KxnM5wPxq4PZypt75ZC6xlEDUldjkg6O+ylYkR8E4Zw7iCFCjb9dzm
G+H0Isy+BqGFhk5JKUwEG4R6B17tjljm+GJWgIV0tdcYtOVAw4jBUcUukmsDPbDhU1BQjLl3LiiS
ZD9mCN+xSr2R76WvkQ4rayW1nfN1A4etU/MTOGhOW/qyoKH/IrTDv2ZqwuC/8ri+eAeSWah7hF1h
VTNhT7ss2+on2f+qYwTGJunbPZpzt6oD72vA0EQ9AdfgIvysxF8RurMqMdHqwVxcaKlNu2nburgv
41AQBibAEcs6vfjMrQMJdie6oEqkvgJtZXyWxhbS5EHmWmSdnd5c1oulgBG4jvCXGPwkAWdUw5nD
0RG44k7mKuSSC8qhi2ette3WlOlx2mbyLbbgztad2NSehvxVoSnusj1eBrG3BIBbm63P4yEwMAaf
p3cFNPcSIUq4pbboo2gTAbaDXfeFU0uv/rhhSTEdR+yZDGfWW4C+TnLPCJtrpBuoLtEj25imcH1O
JD+bV/0PGxDbMhH8Ov8OUCvuMyGGvrAruuoOkDzhYX+CA/LZVY5VTlDhICo47cX3aAFvH65R6sIF
fkN3sVEkDXk8rwDPunS7QzuW0/ZqSbTNAIJQYDaNJPCqAYYPfjt8185ocwPSBOS/K161pXCqIERa
zmoInSsL05JUqc1zNDjTd28zeh6oeFU8RIdiYM9VO8QFfFdLRV+VvbGqTCE20WpAc7iNN42GsOvI
5otGY0AN54u6mfWmX7FLAHMtVMj/abaUP2U3qwkJTIZAQWlzjmaGVkIThNuBvItdgVxUUhHum4/p
iirg5jn6UOzcfL4+4FWLogYSp3RTWjFzldDN/TE/XGEM7WEveXm9gZNDe4srXmYu6xofcNNXEW+H
Tku00wSQig8I0yt+rs+FJiKujwuRm2RiPHfEizAuYNrifgfKV+JnAdfpJF3/GTK5CeON48y5RT6M
MQ40AN/+hhAkg/HFpytKJYNcAu9SIxldnXjgCb4jXE1pCEhIqTaQI9LMK1sxHROgbcblwKOvQXkW
9sIaS/0utvhq3rz8rHQOWQMupOUQ1Kulfsi6DfG3+CpBeTI7QvP4WLhlntQ9jZK56JG54xSFR3el
eXAfGyniZIirJMiHzgG1OLWHg4H5krMNA+B9ueWVk88kRReBvrURRSXfAgh9/mt/6oXWBYDmZ0U1
xwAA+Ism2EaNDll+Icht/r7H5qIfFXxgWJgsi9v0L3iqd9cBTZdji+j5ZMS3BfnMB7tdtog5JEvC
HGINBm++J457B2ErW7uLfDRtxYLqTXLXZDDM1BEzljlFbTAHB4ughGxHT+i3+YLJG37t3SI/G7k5
brUF1ptgWabFXCY96pwzQyUbz84ms9Tg9BYhNrpe6eH0yz+JTfIrSv8skHeIfNMNCV2AZ0d7T4mf
jcSKFlJobashig2U8mFeFatvj0/fw6eLH8xbMsVSWb8VXpbFiqMUz/PEkDgjgMRqf+nONUOq7eWo
7KswLTJI9Si+KFcJkijYSiL+XX33SpkbXVMKWg0H1zCtEjVVz3VbnvBu77XVxX1241W9FnA3BOyr
4L/ck+XBtiOM5ufttzFMFf6lxjSe319jak6GK+uQTnbDpLE+MlGsVjZQWQQ8cu0MdCWOEm69aiHt
izq8gYOfaocQpSeeDpdXXqLv5dRlOBLl+L6g7JAWoFn1Ol8BjoZzZ8M4jpHqM5o8bOX2ziAITsll
yRt+A+4FIFWKSCZjBwhGGZnUKzuC+zTaBYS/lBnB/cZ2gqLyq+ZBti5L7+1MW1uivk18FWvR/GHr
OfelTRnhwXkIngVVL4dy9joqEWkWWOL6jDEvMT8+R00+c2+J+g6Orj4zCwLu5f8iDjhpscOj91fF
7EMaYe4fePCr09Gj4WLRJ3NcJJAwZt0ECSbavq7mkb8+zK7kGXeGBpIEiuion1WKpWWvPVcmtP7R
5gRpng5Eq5lDUJ9s450ylC6bphaH9CeiMqzEkioWgWr6KMqB9StxUlWgUhVrLvTLODKuAmXY0hly
ZoEmZIKA+N3mSurUp84dl/sJWi0ut6SzC4uIKx3+EyK5Jma5cT8JYY86psMQtJg5GTj3zFLoTDHX
x5VX5A0eQIjNQS/iWi48XNEIEahMHluCrpQX3YXJcRlY+b0QI2tn38u1TZIB5E7T7TE7tPJdopqh
4vkwCRNXpMAIX7m5eZSnCKlTCQ/DDRxf7XgGD1FHdvbczXVgYH462TI4XH9Oj5eOViLkJ4Fo7x/N
d0/yeNr/eDWOxfhvnjhR3nLNWz7oDhfQVO281UUJtlqcjmhDT/WOFgZ5VnISWZaR2+tVqav/p00A
wB3nr8hkhLqLxeVdun/RaY2gUjZjUviyqYphRmXk0XMgW/716czQuz6WnEKMFKhGsrufjeSdXFLS
7iuDal3OgIAbxtI7KVOoiUqtnMqb2MwVV7DmqdB0uwu6bCFR1nfpJsOAkHwB+Bvt9MHJvs52SIAO
z65AcwZyDUOKLESpkQhLpQ3DZKRUa9ue71OV7UEzMbXAhpc+COTk8NgXUxuGk0991Dw5NhWKEY/+
gge/3rZ9KCtrv+r2BuogUYkW0rA21qdTKX29SacaRzzif2uINLN4qMiRExIVQuYK+BlwhKc8rW86
nqsjMYN2aYIsvSEBrMK4Bc5ek03tK+9DT2o7pWazENJpBh+PK0haiUVX2zNftTSPotwR8pJKdVb6
tgIy+rmcea4pc6kjDf0c1ry3rImtYGdT1jjfGNCs12IhRxJpQbKP2FvSQCw8tNdrSBUKmFVWkJXR
HaxV2sGT7YXFRuO8/fzuF79TJAyU4QBptCSLcI0Ksxim3p3bHbbDdkpXR+P8P11E4/gyTn10D+BI
t0nVsxfCkDf8uHL2PyFwBdSV3yeU+gT2lKRvNQYt43auaCC++kLl/44em+lSxV415c4XZX7kFUhA
WBw2qn+iQmQ0bcfoxBnlBMTNSNzUsjt0T8Ep3JcYlm0NmAgfho9bLujXSK/NCky92+5TgOqJVRcw
QRFUOdR6RFSlx605jbWL+n8hcf7wCwCMBzHjuHig7vl7HNsdsAvH0kSAjLV2Ikx27ahu/+cu8SJ+
BBRzSD/v+zD/bcaJ/kkGURzl7DJmCXILw6yPdgcOQ9sJgZaoLMpXDqzgmhQw3yHaxp/kAHr0aM6G
bplumlXInJJMue7z9ar4dCvP7xDCODAXntMG44uPfgq+7r4OsiT3dp1WQm5NhiHdSeKkCxYDQhDi
+nxanekKD0LrM/7DcEHxd5sXNjizck5DJs2bNkDh5K2G1I4YETWyL5V009eNNFI9yvh4FS30gUz5
4nlVFD6YRFNKs7+y3BnNXA6svm5g916uG85lM6RpVv2oqlWDdw1wDAwN33wfmORXwnrCDs9r5m/9
HqtEk7ZZSl30unlZHOklZQSiIDoea8sMG2YnT/46P9VFUrSF2Y1wEZC37iKB6VZTrI8vkU2rUd0s
fVf6NVzvovnArckz3DC0xQi2H4maPTZC7MXbYRbTgJm7XqiTaq8BWKp2nER2l9TOFEa63T9VrM/M
VB3yb8Zv5Sx9qOAueLzDXR1s/kpYv1mupkLCY8kxZKF76CsxeFJTCBEwkTCFa0vHzgH9SpULxFjm
QrVRNrEcHF9aHUOY8O5OQk7l5RkLpt6WY2/YFoMmWuAE4VTCmq8tNHovaG7ePd9uAUpCxafdykBB
4s73kzwqMiYhZ/93KKvPMAoIC5ChP02BC6n92ciceQIZpcfqMcBqhcSPGnzHvHBuITfb+4BKH/r6
SsASxdlxP6kJTRAfeDIGmbxD56gTJy7l3BAfY/O8q79gyG9uT7Zpjofo/eKRRZ+0rT94GTlx1mv0
cOv6wFp2S4H8xYz4/5y8QtH6Db2T005mcfJyS5dDEyI+SOITVk++fB3Kh8U9LzU3UohDzn4j8m0R
iTCnzYwkjrbCbpm+vEDKMg0WCKPuU2S5woOwPchjjCcqW8ev2OvS5ppRWhQTCKkRkSW9tJk0KjPl
8FQTCTvYPmRNIPmEe1Skx5u2AJQ/api//L6Eh4a7ghOHWyXjLcgUK6TATqcrNDfifetpUAFaeptO
opXRT6miBsAjrIaCIB71GaINP4F9wV65i+gmrQz5F4Se9aGnsg75idK+XHUC+F3fu0cqxmGVq47N
C52TIHvDAbVdyDtHHrCV46CW3YBg2vPJpH7BEjt/EInrmOgDemB72rXvcd4ZBTX8RkODGCdIdtIL
jcwx1VAS7PyukyMamu4bBIgqYly0poefh1MP+D/fM478OgTR/RPM9AeYrv0HpmkyjBDCk6ir+tkE
IrAnGGlpFp8OFUKzNK6ZHBp1nGleJfGSJ3D8a9CHCPvgI8++CXnYyDInsWrdWEXyNOAAvpsZxnKx
EH2rVrByhDvqBHjHOHgstpaok61wDF+rR/1gOC+LBfvRz9c3e96mlI5rMkoOOnEbdr/yYGG/vJkA
jCqVVzQcHMbZuO022FXPJS6H10Re82dy5p8V2/kuSCx2OHIroc78izskNqUJ6mitmHy628Sky1zE
STfAYkq+ZK1C+Hn122P3YiF9+UTBzrIn3Yo79H7+0ojn8p2I+Qg19xF0gPmSaW/96DjF4FQqgE/H
ezL4TGkKfRp2vYY5pnxp4iFHBC9mtPCnKDzbg7UhXkvsMzHNCvwCiVXWj2QlLd2MV1hDkj8yv15w
wRZVscEoQuJta3c9wQUNWm4iRdpsyVpyHA6cos3Z1rIp1rwFLbY56ZeE9zL0ltBT+WUDPX9Jzj1B
eoX0H9BPygGxx3CoXZWZf3v8i85KQfQNZfiQFHVrvi3aOkuR0H2ABTJIpjdqKpZdg7g3IRteDUG2
4nSYvCYA+y7mdn/qmabgCV+7ffdVTCnDeavuxMNEQ7p+H2trdwNJ8wD/MRq4NG1JvIthio9Pg8Oe
nlgTnTOkB5jNBbuQnR+0O3q9fuqKcBV/yXynv+VQlLkR8LiAkCJKJtGFFD8925zdDCVhDlGgS1lg
G7amZ6OI8DPeABIx6MWGPyGZHfs8fQz2vVk34yVGzWd/XufRZRa9oAreCxTCcgiumWPt+/yS7msG
mEOzITLZY/385X2CSRizIikjg5Cp9FN6hhT9j+vC4Ihi5UL3nW5DUWLiLM3AydGq+JSIewElR0Q9
C0NI4PAxO01MfzuKLQLqcrXxPPZgcoWo60rWHo/LkQZ6FamxhLorVU0ZhMZ/5LYGjecUj8ByI3Rq
//PeX32X5XssUqfJIkzCx3rGDV/oTsmPBY9/1PFcWHVZPx+mH7o1ASv46sVZreepHOVR0oOga5S5
61MvrXkV1IkoNlieMxtJgqrU1eWZhrZinteCtx3EcufWLoviEiUlTNogTWykb3fP7A9my9SVmix5
TgqxTU6gQrHtacfkC5fwNQ+cyrD6ngyuT62fRms+MxYch2Kcy2x5iM2Gy7DloNAEld0bPY3bKaLL
LIZ6nQaYKYH61h1mgK1rsUj1iOLNDC7w3gWsXNgtGtw6NS9n5clm/vhSHbbNkmwxlqsTiXFf/ExO
oXErQSlii+Y+dKD9iGMhVmFTyc8MLZx1nla5OQcLwfy3R0mfi/Kt1s4dACZJymD/mg7uAksbgno7
weR/9JFtdHQspXrEOV8civhI5Z2Q3ivxAywiaWZriGsuBk2PUOomVmVYjih5a/ZqBxttEpv9Og2f
WrcQKlE1e9WpOWz4LWaI2vefFJbeAJGu4VVD6roSUT5lZbiD4xc8TxFBK3bi9Cm2Dr3yS3ddaMgz
bwtqi24dqGsQnEhT+zw2dGvAvlpKhdHDMJd9E6SbJb7l0z828CKX7Qa9P78WLtJDl1w9e8QWCBv1
W9mzeHJ1DMEAnfzGk1fLM+4AejXLb2j25koeDklM2hLvzXkRpcx9Rz/me8vSOw0fLy8js08K/uf8
vQz4YiGZN8hzirS+DREmhZNdeNya+gjpUOuTXdn3B9OmIg6NYobnOor69xdZA2Vii+ZJhMiiPImx
BTSa8SCil462GApOzlUdnD9KA6eXvZaZDtAFJ3aaiF5oX003htXWy4BHbV5cAQv+kuuztG5pnurQ
pT2MM80dx7J/5Di3rDyOFeb21/sPo8qFOH5repuDjaJZ3XyXEHUDDExHZ2V4G+Px9JULN9Bumfjn
WlURwH8fr2yyAsHxZcZrfuZ0bGvIyjW85kBQF/Y1muh2TKWB0KAANvssEbaC67v4D6MBjWyKQyNR
obQXfhGNe4yCJir3RDN6hkpzsCoYZhrUcbeGz1jE2Z3Y7H5jYuj1trdQyCtY7VOxCwOe7A2EwJnH
vdoMmMNtGi+rBefQHomiXmmR/WcdQhOWCkC5dVRv3tx2uuHEQxuxWaswh7aSFzSoz2HZzG/sWQgO
NtR4aXgI/YXbbXXjsQQlzWVIZZ+RoQ8ojeSe2KImegcVS6YF/u3QDP7/metMpzxSBRVMYFxgE1h6
lhD/MX2EURtxhyhwnQV5cET0JZy6yGUAM7yB+Lbj0IVuykO9QirGFFBUZ+xMnlUOKQms6r5UcED+
DAh2cR+e1pRJD64bIpKgscpOcooedyeNTCzu4twGROUwyRHJtTtvh14tFClQAgZqQVajxKXOAkoB
DXdzDLfQYdNwki5BWttlBF+lXiVI7qOBB4BRFfCuc0UuRXqxhOY52zieWEgctx+ZdN7I2jSJ6AP6
Dv6Y/jJjFd+YDJAeHPfWllKrQkL8ClkNHJ7NXColcK+2bOzA0753rLLdu0Mh9xPWRyW0UnX4TmWZ
JPzz7xEdedtpvVv6QXyQwiQmxGso1GKKgl8xPGs904oYd+w4B2SC0nkwi4XDafEyLzVFW53/RI9f
fWVOdrYmpAhmmxcVNgAqb+8YOR9GwQKTvs9pRTMo/PlIDzr06kUS2eJVk4/L12Hix+BieKkiwl8F
f0nnI8hAvuQ1ZkA6D+b5N7cOZ9z8nKjfQJhIjWmpmA3fjS4yjyaypKM/LUyiM8WSxPwHphOL4J8N
VOlJw3q3XgOJ1vjd4mknAY5POPO6aQ0iMAcU1o+qWNM5DOQaStZAZQnGz8Sf9vSuvXDpuzUJAsy2
H2s8AJt1yNEbvyTHfF+93e0IF9H2C7dgwTc9J9xiTfS35cHigz56vBkMWW720xxlrlzmn5Js4eoD
2/8J8IoI1qSQm+fedmx5p5xPZNPdyP8jgnIBPeiXbXeh9Re3Csl6ZvPaLMPsWstm1nWOhbb6Z6ao
E+iyOZ9ZsE4LKNdmY1uzgBV1A54rmOOgqgfUB/rotkSmdU+BmAgxDbpVL+YBAbAHSP9/X5XTFOZl
kvkolas1MTajWXbbmzxRPggzL8+R4dpeHq6173kLeF4pDC0wxq9GmRKEYgdVzkx632eyts9DbX9C
cXbT4NgcdOg6ehpuvMwjW0ExnmSf3+Nnj/iLQplexVudNqW7bFuU45XrE7eJHomNrDXl0Wx+buRp
fI/Qj58b3ttMYk0PXfhHfvss0mCAA4YXiAHnCbS7cUMfSLnMRsG++dVeeS5P7juGFNR7strbbdOb
elSmb94DIt/RsSotb8HBayZcvCLOMs4OT6fBd+OP/tZLNUdmxMFdMdXH/injFqy8rgVcBjhWJoK8
jeX8o6ipstxGw3Pj9bdXks3rHGsRBHGcqCtMgDKXf3IxnJOSp5a25y0cHshixv+Zb15oyqso/HRB
Kkn0pnC2Kzge00d+vfgQo4sVFUBFS8JV7bVCPoKf1IbEHLBEd0bcFi+RXladeCF9kvh6+G4It9b5
f2WpT2iXkf8DQdHrsPGV8UGao5R6G4XD5INeSqsDxztkKWJieeFOTvxdeHr5+DxAw5RVQtoE+kU5
WsfMzpEcDVhEtjARdOC4GMGUiy1j2mpEmHxaEaVZNJWeCQ1/27oW0aUSivAC3EiaBd6OvAzw5Lkj
HGjIY/WY3s1XSNdRZRmI9deyjE7LaXVtd1JLY+NrUYdZ2hhQLfL/zA0NzpA912k4AOL9qXoxMIox
K83gdPkBEW/h5myGrAEWkdrexGmBgRm6eMdRTnZPPP+pzB8DujZobpYAlNTs621/MxO3OXn7PyT2
QW9rBxUEU33FyxQIi+OYFRKqksJnDEfgX9lVMXFxu5Cz8dFOquXRpjp3dJhAWJbbqHlT6djOgUYe
9ivAF1Pfr+zsY7IMXjveVQ8hQuMokocekvpB+kBiDSPa0azTsSyABTRGpEvSoZNcQ+DmwM2LtoiK
AVkj1bRW6s7lJ+eYmssmaV8bI4JMWq4kudQiJJgXu2LaeSj0joMiIE3EE4yPB6ysSb6XNCz2rWWT
bLX7zIdtXowQM7+PflXY00lKLPJPxKzdCYIZlqqNd8S0Wph/O4gqmpkPF04hbd1MqoWs7LnS7lQo
WNLKnIT5XyVAlK9oq5FR84NOrZahYCOSKx5vKX9lnLfHb/MnLp+d0HJDuuUp7t2YFkyYBvFktQ1Z
y6A2rtQrRkKtqYoYejjbq3DJ+38tqKACI8+am2T2xVYVd9pe4hmYxTJSTKH26Gyxm0/9dKV+Xbbb
hTuQp5s4z6ENk4kepqOmGtTk0Kfjk2GvR8IQn9dEdkqlsoYBYboQi6h0iOojSiMn7AQN7QGOGurc
KkICUqHcj2TsJC6TxHuDS5tL41KqzTMCgDe4WkNFODgZztI5uwXzQgdFwEPleTbPCWZCm7xPSVJ2
y/eGyuHBS2z553t6vEmtrbQecjBHKEA6+ONWQQpvRY8pBVx9G33bkLqfQO4pqcyx65sKDzkFwkC3
dGZrnmHXj4afQP9LYC2d4ltkiFcS6reTWCggZ6LCbe1B8KLmW/46IO9OiOrcK4DGfY/6P/4pLCxC
J6vHR3ju5WqWx1S3Ztgl9VLoijNLNHO0EfgyEEm1m/ogbjHn8haIVoCNFwKO+vAPYLjSvVekpxZs
I2A998lUTejW4iT+U61/kqWLjD9ifgLDsFZEYA2xbckwUQXsUEgSi1fCfdyrHsmiaFtefWrhFJA1
XMK5QD9lpQ7SINgAerqAtNL7HElzH5JAqetUjtAYkgHe+/6VzTNudtOA6iB7XzqSu19bw35feEcy
X0HrPIzb8mqhphKEy/jAvnB+qzwUfQQkIgxV/cmOPwz1nG6Y6Kp2Mnv7CewVNIM6sbs93VhiiEZO
eG+sX/OY7na6VEF0I97FjhTCTNYcuqpPLDxxE2DLymEUkswLEUz1YO3UuWOLTaXWNUgTNjRLpvte
mH/PA5r75Eao+B/ZJFBTrEguzcO/6GfZvROBJAatvqr/YIWuvbaGFk91IgN1imRwpS65Aptzyu7a
kWjT2/XgZCLzaJP5Nj59VxloQC5R9lrOenVQTsqDJzaCHzAWdifutaXWMpb76OZGs2KjvCBtzWhq
aYmx3r3LU+z4FqomLegyd9syN/nBuDWA//Lm9VSV4ISIspFLxdOuahgUbUn1df1MZK5BDB0v3SQB
wylvjjLKqxIxV7FATmiO2qgizuU/uVLPtlzmO4WCA8ZlC7ZSMcZbQsQQ9fS4fICWRrhJ6hZZ5YjU
VMHvFOvnrs2HAQU/lu0O/W6kYdKlklRVNq+uZXLloVZKeRUaevcgceb8+L+JYoVY73gYZHBM85eE
vq7SZE+qIBB2mdzpFkd7g1XUgZwrYKmZGjvJ3txsUYFLXILIiwS4DkaG5sG4AWaiqnq3xSdKScch
WaQMRESD5vkBGUG5C3ANkvpxsr/JXfMScir5u408TJJNQRcjMWpRnXW7NhC+dFgqz9pKGcTlaPdD
zdJcrZpR12rLDFE/L8xkHvvhgQBSoFPTZRs9mC/1Bh6oJ9nvSFOjaLtC3ziUeEBsoqY6oIliQ5Cg
1E+r+HzVQeKiDwrUaDVR+91JQQ5UspsiwPJ4oza7Ws/3KWcZgC5zfEHZXTF9+x9PK50LXmfwLOdV
XHq16xp+LkVjJcC7K0Wlj3xViaXyjnwXY+5+MNttOLggS2kxKcGdcUTQ//E5hc/CObAbMK0o0dHR
8CtMV6S6S6nPTzMoFO2URieDAxV3lZGPep+7RsFTmjuHZ2kvWAkR7dQi5nLXPSZSi3t8CDDpIVQa
Erl9Ah9xEESK0R01sMC3tyKm4w+VZy4+3ImP6hyieRwre9D7AAUXKXqn4HWrOSkGjgyikUnE00Iw
pMPUq/mwGN2tU5RL9/hpITceHWChue+1DOkdW7tSLZcptkrAM6DnUxFlkRYHwW3b22LVPSd+EeMr
n6GJ4fkhVBAFcHVK76ojxav8552uKeHhjjGxPauKbEUWKV4FErhtdpttI4L+Z3cED4NQyYNNJhR5
tP4Go1qO2Hf5saukrBp210bTMI8wptMr/uJLeWlqP5voNv+/1Hffsjh4dlspmqXcoBphGLopa8vR
JTQCgMQ32dBScvpyA0u693bgMuqd7Cdd1ia6625+JZ5xEznHswr/hsqNSya45/bF9rZkBGqY0j9E
Kfm0AhcOCpA00TwRS3LRVMyl2qAMemR6wb47mAi5oYx4+1VrIq1vRQxKLZdG32B/9iFt9q3uWzAF
t+nhiO1I7Pb8ZruIDNvPPhEHOBH1478D4ITCmrTrlmKVIvGwZ3AGu4UIuPhigNlBoL7lCG2Hn+Di
bQ64MaAH9d9wmkJUWcmiqabHsjRAMw0Th6idoDVCPSif5WcyKGmMA0VDpZcOCv79dgkwvuzsnSnP
vMjlKLoSRrqy6WuCU7i7n7SfomLx+6SM8jLSkclLY3f/OHHcfqSZybGHRPZwIh70vLgB6Fa0AvJL
IS8hrhceQdTGKK6RQ6R/qIlgoM1cumqj8ssnYLiokVfbNRz5Mx5fEib0ofxqghp1/K6MeUONfhzq
wqGMOWlo4XFQFqm6cR/N3EEGuqa+mo9881JDNXx5IykARmzLEBQC882FPDrnQbuR+3PlmYgDb18d
IvJq9lpY7z9eZo2NkhH8l3RQmvyG6ATWI1RxMiDzAZ1p0OYrtQnycurCvcT9A4Z6AmXDZxZ9zLBS
DTBi61GGgdN2UZK5XHcg7vMFATXPKoCU+Fv6uUl+Me7qnYHhkd6PNMh0bdq/7kS7T9IXJMfNfmUa
dAYQ9YJvivqzNW6Zqk8RwrX5wvV0Im1ROGKG/u4ZWwlcwRPfE2oprEYL3MpMrpQ9237lAR3p6X91
gYL7vEpWvrtnlp3cAx6xSYKCxfz4fUt7ZnbjfYyFJhy+v2FXE3Rv9NSkwiK23JuupiIuMf53iJEE
iqYm+gi6Vr+266SD9j9qSYkV/rkZtYAJYL1IVeW3KfWWStUvhEsPn6SA24QgwMpE+2Iy3YtGUKnG
dqPqGYhdES8oKzGu6Jx+PXSh4Xy5ew6UxG1UZb6+cWiONz5P26ybGLsaZQayDCtYOhrcizgeMban
RAcOgyDBk/JNbhz2tqsyVbHhTqJrDLWQC++zNtBFZsOVJYQJc5jQtxwEnwOVF83ozUNEs8RVcuZO
FVfiOFUlnxH9SG74K6jUOsaKEULGIGX7qCH/Eo5ail2LpTf4g/qJ7LWxURavLySlcLtwT7SGjccO
e3KsNKX2WL6UuNXcQWUREbrpA1zrCoO55MNx1IxrRVr36XcnkuL1Ky7i1M2ZtUbNxzInt633r+ke
1NYPlmbhFfnusDLCzolfoZL67zHDiBGDwnpncoAyZmfcLfWwUAbp2Uz43MZixQVjTHZmx5RagEz5
wJvSpW1zGQwnL2cZCkIl/eJ4raJ9osp63Y6EY/kyDA0rr2/GLZObYxegNcqGdM8sMAtsVoGFLBSY
iVx9BMIEUJStJW/jFCgg5gBr0DMz2bFY3aYvYm7VJN1nZewrvuC9BSnyU7pbGY6S04wPR9X4XCq+
vKqY2afzmtV/9X53xvXCJGSyq30usjwJ23CFRwef0GiLg+6oAtQG+j8KWNcakVsUY2LDUwPys5xm
EZsn1iesPXesgV8SmjaNDVHS4y2931ISssWcB/KdmbFIQu5VDlbC54JANXHZitWueGzHV8yqCERW
ND7u6HyFsW1/90+ztxFAHH+pYE6hdNNZFv/8GatNHCJi8wI3L4HkxjBH7ZABeF8nPzRlAGiT1asY
wYm9+8H4h49oWHNMDdEeRW5gwbCIEQkXZFXGblBsNEokDOtbaDy2u7adEOEz+iK11r0EV4x27guN
zVf7okFvPqKuDNRJ7cYa+F1igf4J97/Mu1+ACSq/LaWC6KczDKZsQVlgQbX2URUK3/+18dv0z6sP
1UklwnoR8Za/a9wvG4qoYxqLXmXGZdjX7/pB+Fkut4JusaI5VgJdfW/AVvF3HWJXRfvzamKls8v2
xPMCtoHBIWD+G1504ptgiWKPCNxh/ASZuyNrZyLD0hc9WHUcLSFbu1RFCISkKAAtQuzD0KDluPl8
cdJaiN8pZBMHK12OcejSiTTwDLiQtenUU0Ulr93tc+P/cGinwvPHw9RGQYgJ0kMZuqv4Zk4gqbwa
gy48gBL+om0m5jjIGeAbWdwPudEalhBIkgchaWg26wCGzE+782C1O9eZrEvD4w1l41Td0xMOp5ZC
TlzyRyiJEDaFXyV/YWqwNy4yKQueN/yg3RbIhmnRJwIcLxQZIWJgDxQmmpcPfFf9ZPLcBwBgT+Im
7g5DvK4+RNH+FBSgjANwRHp7FD3+Q7FkygJ7JRFnKHtawLdt64GGZqp7MdIFqjpgpJ42Y8cjj/1N
PYPHxgtwQCR7I8tebZ5Yz6GYYAp5kxhPOup2YdPyAwparotZ4D74NyDMbKRGPn6OG2eKZbLXsfgX
NHvb56q7F+ZM9vfNcYGU4bFr37bDAJM44bamrpoYLHf6CZ+/+Bt80Y/o0+vnZNG6p0hxqBGgn3Vg
Ov9vNlLFvuIfrxqPeMXFewFvdePDEqN366Zct4rNvvKnEmlPuCFKrbh+AxXWed0IsEAb11Bcvddv
CCYMaoWNAa2SpyErMQPCO8tuxMVPDk8zaMigcCwjeqM8QiVmBu/t7gxJBCf8ovqS+Is89rvN7eLQ
B2145I+hcgVe/UxQhJKvYyGQk0YNrY3Sh1VfA/KC8bydW0qJLm33hq3unDuMkqz8sh2pJ8NM5iO1
UWRZ/0yJu2lnDdlVKKuAzGw/m3INGQQZnCo4x1IzVKsI4rWpcno7aZhuB4aj6PGFFc30edTd9aB+
xVNExgC2Oe2JqGnLtZ2BqOxPb/8/uNko8CD3BXHCVgqX1vR8mN2Kiv/F5q0cqMnOfR7R3KcwLEI+
Mvp9Waycm2MXIQiyDoNaRMg6pGC/1esd6MLcDR3UyrJWJSMqQtpkm6hWB3fCnzOUA1c3agfRBzsz
AjMpBNV6RA7d46lDova2BmMIQ6ncqMtX0Z1g08AFDTMuSQM5y+V/PYNMovGzGZk9kJf0JPLBfFOw
M/y9pBn51NSYfwDzTWhQ0ecm5sUhGlDR4GkBct47xfTmanFDOscrhwsZaao9L4G9GzSWs915N/ir
kI8y/J2D+9de+/c1CupQUsbRDeSJC0DdhO/l7XadGqgUrkA9FWM8MBeq6OjF0L8MJIdqQ3/5+cwQ
3aRKFco7EtUaYIVNkRX/dtOV3uqz52GBajC8WiO0kybHWwBtRWh1thZiJTXG0rq1lRjwxpmrnWiu
ACwxp4PIUyYg5/SQKm7rMV2S5VUD1HTuI/i4EqrFwB+mbFvLKBRGRo0yw42kiX6UqpQ45IgRTIrP
42wizi/eNwQmdnB4Hzbl7cogS98d3699p9/pVCE3+nXQ4Ho1oPxb55LqOvx8AlP5yxrqQTdsdBz3
jmFMUJLdK6Y1nC9razRwtnt36IoAABeatRtJY5qDVbYoyPdCa1X3giq/qBg/hLm5Xd/LFESnuuNH
embvxOFY6a3opy5aSo2yCvohA5xPjvbbK9tz/F3wVu9rr5xsTr8W4koB6jZ5c7HSRnuyYr4YId+H
TQUXqzerliJ7OZxG4YYy8YxH/BMWLVa2A7VYxxSHcL/ffRv1vZIdPQOD3W6V4CfqbkXV0fmbgViP
Z8TVRjgVeMXZBuPqFGDDgcspNItks3Tbny/TB50VLcAkqyHKwaVWTxHlUCDctOT4IgkYMD/wq6+d
P3wVIirR647Yiwc7QhKDRzrEYdz7fu9lccjfX83EGVI1LjPL3gftG+W7Vqf0OFr88ipl+iE2ACyp
O0vUV9rGur8lcd8m0eZDUAlMC1YTzq7qc/qbwdonU9G23eNNpk7TfkGEgL7EjNY1F7TDc2cDZ/UH
u0yOrhk9R5MtLHlxZM4uXj7pJHnWHOtDHG/VQy5+pfow1aTppsZpiM0yq/B8zWrvCsym4V5KY8Zo
U+0aDt3wp6KAhZSiWsQe1fXBLg9HVsiO7MkGXVKMnuhy0T6qbWgR4JvvWrv65oSOgISkajdexNBY
iamI3Bvtf9vBbRChVP5RyOoQL+uH6gnN12Y/d8V8+x+PuYzQbnTS7xzt61/aTm6E/p9d+gXhVLvd
heULHb42xwj9NyoyJrLbsJdSVs8uaffjsO/+lw2aJGgRT159Sm8uRIaBPGFuFECmQgg084FKkJIX
ae6VyL5yN95xoet/vF8XkqTOvIMRpsReahmGwEgagIGFiDaCYNq6+whgwmejVoatMN0eTFqqMNM1
0B/ovAeU7RRClJJv8pc8jj0tOlj3jyC0pcPxODQPe0n/NggWi90OU4cxD1VK1dSvV1FvZy91azDk
ZKFki7WpV8BjHo6bqXyJrYdYdahlb4vudQw+tPc05Zeo52uD8EL2ctlKWbI/r2c773tgiHwCHbF7
ioM4XggGfPYQzbNQP7BUhcsraWOmHfv4PpK/a4XLhT48B58RAEPGQaCUDOelEi5K6QFQAf5l4pj6
O0jADq3y8nDpuLYHnH2x7uIgxWdIzMRn91goxZX2lZHNPb6YAjRwCcS+q6/NVKXET2A/aymk89eO
UD1kfgcki5d/oi1t9vrkM+DVXph0bHxGl7/4JTuXyt05PCMXiHcQ8mEBoYNJuBQ7PWDewpFfRtYu
WFibfF2kJCgZ9+2gibtmDy40JYUpalPGRG5PRVYxsP2tI7aH6biv0F0yAaZssnlK1HlIFg2myyRF
6mFkjH1qsIirtObw5RK8XbT/gYI8F5E6PPMXODsRXcKnpZvuBIH34at+a0Tf/9fo6ykE6PB3adVO
0O+qcAsMuf+IYjbVIvgJVUvY0F3kPEWJnHzfBuhlUPzAcKTjrq/ommEoQN1gvWVzC/9WyCI3wByz
Rp6C1xeIzQD45iHaQR0lz6a4a3Mmfc7k5ETFigfaS2fnXsqgaljzO9d+9i2Oejjqfhk8KuEhaizR
HX5E8sRzEhtDoee5f4dDCVgm/shSTz5rXTYRLsujxCK5ZR6jAexHzuKrSCW+GhXL66EcYEjgNPxW
oF3xJTNi7Pv4tqzhSyLUNVE96Ndre2lQ5aQDm/WLBwYhMYOXvbOYkLvmNBai/zv/EXYAbPtjgTNJ
cy42tNu1pzYeDsbODgBvDtIeDoPCHMx+wjxpZbdkTPEappJj5VPVKAoLwglgaroMjD1SFdxLQO0h
mK4uvZjEQb2ANbZD8v69Q6dc8AHIH6ZEWUsUJJP8mR8YSk/r7Hjo9h1YsMAgn1LfHNgJGN/L53uw
w4w13IV8oXiDAekkQpUrUWqvkpH4CAizzbvjacL2+GYT4j+sxlW1dk3Z6c9fsVVGFwS/oz6BGnrt
ZIJg0pmIZ1BynNG8v/BJajfwTkC5V3DUDjlErMmvzuBffDDMN420aj+UV4fMEvDwnKqr/imsc5xT
1jWavxy2Wmt+Oi4Iz45zpeS8OpTI414G71BgCjK5tm0GkIfAJBSuoBX5OO8LdFv6+Yrn+hIjTNzQ
2nHvMbITerFPBA/M2qfCCi0ItaCHxoPqzOFzKFxlOQZvmAiJ65dSyI1snHx2dCM7onBShnwfM25S
GiEvgbxnhwGGB4/9HVBzPEma2ooHfBvFhnTA5sj5/6+StY7hymrw66vU4wAMurOJaFuL0+n2Y1XM
CB8wn/7w9fS9Lm+m3H6WrL+J6pondoGkwDO4owp2uBJvAnQnaDwxRmTWXaYoEj5jYBGY9Gw0zY3E
X5C7KAORCdhtQVYWlp2GK2VqORzBKDTzKFjp+jc4YsKt5MQLfGm/abIYXQlVCzhCC3vFO2b+le2/
6v7+38zWDBcMntsbNRrvIwScP9VVX8ArwsZNUqGelBQALwZQTsD5LI8N6LwTgnoSs5qmobkWnjwL
bfYPCox/dwYKEHUgMxR/8V57cZ+4RfjbPSMptZuk1ZP/v/uMa8mk7XiQuE3tt1dIayNRmNTW1VwH
4xe9aEKSVcCWAxhMCiBUVxoFzuwySAzbCuvS5sKAGt2ZV9x5t28/KOo7gBuo1JmN4ocpSsYJGPqi
25dYDnbERi+/LZXjR8OVCx6rZxC4yvKCC8Bj14PzJQ2n0Vzr6Sg7PwEJ0r6tXjxq8QD3MEKdytnV
Muqyg+aRqiksOO+OyVpHWLBvCCfmDnSbDtChO7ZV72uM0AUMvTqKK2HEIXMYtLtssKDlT0Vx7EvT
re6R2QvhkVAJlHaB7aQcJR9Xc7Lu70ffnWELcDWwR5jK10iF+oI293C2J5845D4ceMITH885+ZKk
U7e12wN5gwwrFXe0yvHsE+lZU6lUKzyEdi2nMI3yyVc1/mNa5qm+hvMMBjKTy28q3RN6HHKp3A96
FFc7WkEa1Bhj6QHakdVK1DjyegwsqqlDyBqtwNv9mhDbZ1MkPyuvJMQoIHvfNSawZHfN3IBZfbRS
k7YC53k+jSBWjDkzOLGv/B4SH5NNBHwmhyv81Pra8MSH+ePdmmuiDJKFG+d0nlvD9lrO2Wnhpvxh
zFq2jBq2XK5dtVCJaymBbLgmZMfZVxjBjnpPXQEN0QxxUts/zm4c3iWGw2HkAfOeQe0Sf05gD7uk
mRo3Y/sfEwaxVit3XGz2Ebu1dKkEm9qsmLvMAk/5oQLx7k0hI8sgdHT6HGuVdZB3fDTd0QcdklA0
/GVu/mfAQHDZYR6DpFxn6rk8/Yi1SVykDKHqw8WMAkyOoO/DIO/FmHO9yMvi1+SodRfh1s+YmMYj
KHnxfrPTWaJ6FW3oYaK23O0BHF0gAv0rmE1L0nVt7m6H+3pdr6PQJZdL7x5C7DlESDzTFtmKHyUW
+5fK8Juq9ZI4mqWaG4wjwbFtavtBVxwPczFXO5brzaiv33Kx2W4oFDEFR5oVLzEXNlh/5L4IPKjZ
Smoc6FYszD7Jc9hQHOJYl/XV40CqsWDkbvuDOTqrKzPDkaVRruu1++nOew5RH9PSaaLTCepXOGLG
jTuQHpzvTeO2BkeID7vChZ+4n4HWWQ6yjLnrePS8UkbIafEHL2ejiB24GgENgfisI3lwjM9E5Kga
o2uxK1f5HtkvqzcvyVFseu3PPXKWdZKoaPQLwbqs94jOPDVgx8VLlc3GnP11jQRB3iJ5N5igrqVH
+L/UvLjet1xV/HvZJEguhfuppPBRoTNrdFeiai1wnM+vYLKmcT8NGJL9iZg1PrBI/LIZLT0kWiqk
DstAEYVPD+nWYQmbbxTePwS6liCRz9iT0XSydyAnn8MxTn+iBLkiMq7U+HesN6P8nLNwulwBdohS
sS0vaQRnppZhRgIUB4Ej7mS3MeBAPnzNWsoDgd3iRi2bVmCqff8tgom/1nhAkLv5bPvDFPe4Yvzy
s8r5/qAZI8H6l4mF6h3QJ9uFdrQbo0XYfd7kjd5B6ASKeZDKobrrkm1vj0cvgIxUOyjkyptihYOt
h2RsnshE3o0OnR82bAW9AO62jXhr0B+uBHAym9OVFYKdP81Ek9+HxdUNODo0KKN396jXjmydCHZB
Uj7o5uVA9I+ojhH7rW5TrYkEzY9YWUAKYkPzVh69e+VRMs8+SH2D8Zgfj7aInQbHqO6rqwE+pup4
pmG8Q9pF4a1PL8cgWd8YzwyrLodLxnpON2xnAysXZ9Qh+f+dIdO1TQHjTBa/TbNgnKGnNs26KQ42
8bykwd4vs34Z4kszJUZt1IIqjjUDkythA2IxnDOaq//MFkFwEMHJynbiOmQtFsjDXvZJZjhxHFcY
urg0HOgPBEfT+i1maPznB5BI4DoZWGGvubItxK9O4dy3qjzEMtfrcLWFz13d/+vL2whZF8RYbIWI
yGODhW5RmHY8/0fUVRbEicjtRDPeF5wDrJP8bYNTh4mGDjH5R3x4eEy1WiGBg6ziHxMIU7Y3pgk0
DuKhS+08cbZxmolRWbjbPFx3yarBce5maCBRtutp1v/1dY0pJtEpHsn5rV2m9e+Kox02ZVS2LTjo
Tl//AD9cae40mPw7AyiCM0GE1UmppkvVfXntuVnW7M5DIqctMI01Fx6CPI5rsbx7s9orr0eNhJd7
huKTV66yVQAD2pksKOlPlUsgEQPbDJkFHJwMJPCIUNB/KQMJ3/TYI30fRJT08CtDm2PiY0ORMPWW
GNEgmW2VFGpqasLKjdrdC7x+WjwEkNW5PK28ZkKNDCqzRY4jPl7YZojh/qcqWBjjahjaHKacK+rg
wjOvu7k2MRMWP8z+dsTHaAE3Y0Ggm/08l58+lDToac6sZiK8iQlaMIJOfmgLDIrW7nGYKvyCuZin
5dbxQZ8HGF2qiagqon0b2pxm6AW05zqYYsoExwaL32plYzwPxksJP43ewZzMAQlLRJeGS2uzwn6m
F070gxII4JHXLXQVRamtJFm1A6IvBgCG29kDJ0jhglZkEIGj8FkbFRYdvtr00cmbx1Hrael3GwVr
yu1bDyV0SsM/P6jA5+WcrWgVpm+ALzWIxaW5RlkeW+tCcuq8wgo9t0VSrEWiykDMsJU48WB4ssce
EmMvpK23yfLR98HcyYKgDLgWFhSRROqRZstN2OxQshDrJZyA9s2wqf97uU7NneHVPp2BOKpXTMAY
EnPoDgYzUhneK9JMuR7J7/BGfnxFrcIazWCXFOgIpAXnoMDOa1uXLnOc0mScNEDlBnM/LrfQlMao
4KRhUNBf0o2lnm28y02WtauO8NIYb7vxyBEB0Pv60JUSt3YvlLR2JDhhpYagLK80A+NKP/ILaZAc
OZCRG5bxVWf73De4MjQcXhY+y8mWZd9qXXsM/mu4Ep0S9UjfV1/K+RlydwusSqrXB7PiLoETVw7U
72n9gp11O905GUmP19b98N4agqyT0MCNMSPneLHYXLwAorzdOq8eONVsK/6VgDV51WvvBDgtFcis
OjqrfQFdlaUm0ks/XDiySXDhx/KFGDf7BMri589oth0Ut58MyllkWjN/XkX7G5eN0DCL6Y5tQkl2
WjZW05wgf1nm1e+69Me1PBkB4FEE4MyzndmL3C/xK9Wg2lkXupKh6e4kVQleXU/MEd1ozAhoHO+w
HHc4Y/+zbgyKnB1TRulX/6otVIFDvtIrEaLFjMOfNxfI2NRoNnCcqwcVMZXkwuqBDONtShvviaNO
tGtDWEcckylbK3FucrD1k9/+ZQ7JcrQyI5k4zAeyNyygtubMjriqsBvVIRAVT9r3r5P2rM1ZMOAs
x0gdx2TPBvoH0CQMQwz3FrPftEpS0J814/MrxrWOzqUSAFriywKbdSE+dGF8b5baV1657O7180fX
msZlFOevJtxa9TF99bk7pxCRimFyYBl4dKoPMi/YpKzpr/jS2yfsHLgj4eCeRMmhoi0OFpqNGqWG
CsDeovoMSOpQqOV4SEB/vpJRjs624X7sf2Q0NZZ2olkUIXCsKr+vPETlQMLf8Xytc8QRaN01RVhK
VBeTZZSvQn4q7A4H3VCLYOeaod27cQgfMhKdWOHEcYQJBFGI9bPzonda49ZNPxMmDGzXCdGZ/Tw4
34Z1vM2lGAoCyTDM2HOQSqxjYmTZLhdsdlL0+/5BnbalPT+dqVYdu4MllcIjSVkvTX7hqHT11n6Z
paihIGML1IUsA/3CcAIkQ+j7boRvKsbW4PQQJPaaK9g80vxnEmxzrbVtiZe5+kyCrir8qmjU/zq+
kXvYm/ecLWiXHqcLw8XcPhnaVR99Ol3/XybRroJ0HxA2UYPwqszJ08VhpWRKMZbnqRHBbe2fABLs
sbl8q3O2unVbS+kkM1/jn721VH2lArfEeSjoVzLuFIS7NgIeMHmWHA1VOHUXFhIudGaJjStd3fny
TuaREwdWNbfm4ixeQ4BfAkDSy42QphdZiNnXY8XcIH2ukBjPZ5injjIBSo9dqmj0MzSbCvlCAtF6
Agp5oyRZOrgHk1cLRIspIfzxgy/McfIJZIrRvv2ySkpfPPD3W+kCUYqLZ9TZvns+K1JCafEpPdvQ
eBxsLxtZs9c2SRB7mjVFoRwypZphlq3mLUF+j4sPXfvYO8S6IDFKjo1lngVRXC25Dr86mwGNv6z2
RJtiSHPNX6MPjQN76pileW87JVTZlziylFXTwybbCNAFgYz/MWHJJLJ4nvFrQmL7Qc/+6idFRxGH
SUatFd78FtHXes3bCs48fJG/IVQ+9Spw2EyFgcomlBcWI7VSyhfrH9SmjAn4vAl3+WBCfFwv+jML
wzEfSzTsMad0XKzMjgsztD9fxsDUMGtxmeyrLmVnPN+re4D0uIL3KfnyB7eVmLhHJLpJUCu0tk+z
cFxfjy6EUdUd+kuoSh2J08mteON0yHtys9S9Z+9gVCDj7APe/0uY0pkxurDyoHfbkigIng8gRGJW
yGEOULi9zMl5HZ3HLBQvM3eo2eGmyJJidtXkNkpxt25y7q2v+U3Y+0tTkDt60LEuO2yRDeSJbTDT
oRVgbVmrFx5azjuko6GU6mJOjzrGDP3BBgSjdvwrZfjT1lf8AjQAlgQGZU1oP/QnON+8GHlCB38V
jopSciORLtwbIIJxjtf6IPhMWuBCTric95N3T6DqXIUxsFmnyNa0yBdnvuACPe/ZqP8eq5fnM5vx
h1oBAe7gagFIClU3+yo4apTptseNTHhgn5bd8mwGn00HRqe/bu5RBIwEK5DnXGLvr8fFZ/VMrhiF
chlL4XZJDVdJq7VKwcP3hNR4cXiC5Noll/Roqb5G+sOvR0w1sqijxUAHx+JoyWEnM2F+VTmH2lAt
isEImWrzEet+1rOjN2x+6XcQbicSFaZHvJS4VYLqKbUYueohuaX6Bm9AFNd367TaSt/Y+r3dBwoJ
TPDq5jp249ChIWdNyGZTDfInUNN+IR/HzCbqXBuUb+jtr/TKMSiACFpaKcjkKgAULX0SnAtClIXt
KmqOndU1GMYHeg3IXfhoAxulYxQCESmGUwqWQck95Y3YDiZX5r0eonrOaeACE/bgYmaWhHmvWXaA
oNermzypeoKLZHxWmTRktu0wpT9wNE0JVWv/WkBhlMXtGc5w/pSpdj+1nnJFwDmcVBnjav7sEIH5
tjVrXzNGt2lOlAn2Sl/AmuTS/jD4lEpIb/KIClSHqG6mfADDthVBV8sNBjE7iMx/YGKehIC04Zq+
gqgIprPdBJvb1snAly+tSGA+PCr2GM+HhPUogHSfftWXJKKSUCPtMTn/FxVrDHbfAUux30GI4Z9w
hoH268MTRcq2gurhkDIGG2XwYDDM1b+IABSHNTdpVcmFTI72En7f0wv76cd+RoT1XuyqJnQ0lXRJ
5gO9UkzP5T0ghNr47//K9+0DMha0zDBvn8ePZgMxreDl3VdySIcvqU7kCetJkyXqZ8da7JBvoRou
SB3Gxu9IjtKOpA4SjGXi2UVc08uSTbnq8S3LVWpXcJmGiNona5luXomlG56jgX7y9eqYauy/xrIP
6jz2nuu3GHxTcADDMTemd5MYn5NWsnrj+JaPg8JRqpUnAVTRndrBelDifj7JAsLZDySyroUoAqOi
Lsu/Ol1dEB3LPJWtLp91+AJIuf/n+G2P8WL8p81t/9cxWCd3nq2N/Il07rLvdt33i8pysfVQIQEh
j8zicZ2dw6M/kK6QE5saG4GrLhJKxF3fGu3JxB7Iafv6bpZxKRH+6X0aidIa7j3KW47nvajwDpy2
4TWEToPsiVuoQwZ8UvMgQgI/0KHwjWhf6fcRu3dgQ0+nrVcMG4MBybRmC4IVBB3AMx1um1FNFCUc
d/LlMzlc7xpZi4NY1TnM1xXARWKa43ayYv675q9DHdW4TqJvzTIASBl81zYs5hHc3XGwJ1SsUu9E
2z6zUFV/fuM+2utJK81RWmV6U9XSmnxRNLC0N5DmPiuGyUnTSaVavVMzs4GBHmYsXHNl834sd7cH
cAfxmxeseNF3Ohl2ekzQYcrtHCjuTeUCh4AObUFTS9daKK8sc7D+ov++qrwPhfBMMvnkUqgRVNg7
025ockj16xnCnmTlhjQGp0lraldfP3H0cLOJOfNIepNZlqyV7m7vtbdtVnUPYEhIQQ09FCQUNFd6
cab8cvV/ZSf3x65NnJNtrXeSu9xNBvx4Wug3v288mhiFRpnj3EB0Si+2dL4lH9pFYSUKUYrLd3QW
seC+533MVHwtu+yquah/dbEvYridtc3DqLyOmKXDMbJXJuZHHBHRx8bxvsuRzXzk+fpLiPxv3qka
Ozp/CnxXQWjiSJsURGCP4xqS+QwNquwYeLcdseNylo/3/zOvTE6mQuvnXVgdN+fDdelQ0IS8jyAo
0Uy1F0M324v5rtyEzxu5ZgHPOIiQMRGruhLxp0A9HCvh8GCLHbdhPq3FgCCGFVmLKzJ45L6RrTnw
Wdmzfl0QbYkSGUbBRY16zxy01K4AU7vEi7ESKvGwqYDvHYRvxkUgFkMR5ObqRIcMUmytP15l9Mx9
ToEl3uJCvRomKDj34hBpt+7PlYCRGkzara/pAgcCDdlFEf/8FPNGxVXepqgKU3hXxqvM5tdrQRyR
9L1V9fGbH/g9FjCes1OPgfFbUEhuVuujEi0rtG5l6trbS3qJW3M6V23GA6BGUMMwv4fiWMCsxVF1
UuUWaRmUNoBdwJU1t1xVtGy5RoBOS1tFHsDQvzs8iS/B6d4ZI9EQLQsYOGysVmDxJXDWserOQib1
Q9V9bAAE/0te1eN5FhHLW5VyfFsZE1O2k61BeCeWlA3ugUYnCeWoIxJXH2QVXvZ6C/Inj17wWvuD
e4o2IQ56xSzGtaCJ7zT/bDMlfFm7CeZXBr4C7EDr5qGEm8EzEFZ19k/20Ua/1+877XepcepaElrl
4+I2hM6GqdF3fPqQFfg1hswL5mBHdPj1hBppXkDwocXweD+Iw/bdiTxzR/pOC6QWZaeqPz6rC8w4
6luyOrCv7InLic2qhM0W+n8+4aVT2L+qD7v4aMN+BeR+goyTueE/dQYmg9cs1jb8sBeHcvdcxggR
B7vYA66RMiGbmjQltuJLIYtOfRnsWQW9gpok7SqtuYjP2D+O2SJkZWv2A9w0ITNx2Ti7QXq8ZnBT
nPvLCgJHH4iMkB3DNT3/AHZWHBLSB+Sd7bFzgQgmD7AnMJnS8LIAuOFnngHpY3+uu1ZYzbzCDjBY
yVB3QpLTzZfrocyBalf76ighs32Kyoph8UmKYWX3mrPRl4zfqQQw8iMDyD5e8ERoUZ2W50496tA9
vUDwQ2IiCXUufrscxUC/iKy/AddOxc3x4HwMsD+KLoySUS4S6DkWangH32pupibwYkjqqNh/Zv1g
wkl5aeGXWUG5q33RuGZSI/L7EwYmXMGT7776eQWZMr7NNfjudH1DjpVOZdpuv2mcz3dgiABZAZ2a
WIc4Nunw4ut+cpQpwkHp/QH+lEPHOm0fUm/etuyO36yI9cSMZms3tgVvMB+apzcne6BX0Q2f7Vzv
A9QuLkvCxZVOCM4zTN8zk+lBs9asWGU5+JLWSAJz1hnJ3Ri1Pd+lpVncNWYprlmJfH+hJueiOSZH
0XrZhnl+R5Zg1N3zjfRAovumUnKSeLT4fOhE1AvOJFl4jp279cMyNDdzzGv0ox1maByv4r/9f9Mq
Wdpl9mFyla2ZfJEhRx4YZIoNeS3gBvRYfRdV+AnN14LcuK9SsxkwGVpLqHprujJXfJlR1zjBSWs9
CN1+rOHWzAlUOelk2pBtn2oHFyeCbKfYi8z4d76uRvHwgER2fjkcs6ApFzojNH1D2gNjCaYJQWd1
WAWa1QI3cV4frRV3o7m96lzfcAF3XlXsWGs7Xss4e5CE8sYqMNF6yH2VNJS7oaae3G1lnB8iyQGR
Qjg9HddA2zZfwaaUWi0m3cZ+vr15dNGsnr/Yxm6XlbSZSuVDd1GR79PnmUqdrJQhtyA4p9ZXCaz+
GpmOin5g/TnTn4WqzBvW/4mDtOfAe8ZSitFgjxDEjFk77Mem0QnK79JFmJ3p73vXqlDY0ZK3K9Xi
Ryke25NLGCJSccitguYyTS2iCKTCgIqpKVOs0a4yatzrZpvuer/jxAGhlNw8Kb7iVTojegdrkl1s
UmhNXyRDPJ86Wm3SFvy4SKxQWFM1t+julEIeGdAI0SDo5VwmXDpfYV0SovzJwfNRJdsDOZHLWgnl
1HlbI1BcfRxqmZUoT5jclsUupTh7KEEL0/jEPYW3hplAOQbVc613xhIMNxQ1nN4jJ6NklH8R0WpR
ZEMc20HiTBMic6ATvZ21HnlAmJz1T2VD2EtKtz7LFkE6RbpUv75xp4EuSPV6zPolNxB7A+uMygeR
RtFS31jplMcPlUXCzRC0Z5k1D8Df4yw9x8SORk9NhYHgqI6gBZUpIyOfo29FKfohske/scrWcS9L
28fsQ7gbBujEO00tfOrhUwQQAOfZtFP69WpuJWhRlXr92IXC5eHMzEc4cKHKimv2IgInbuXAX6DA
pplaQAVvxQtNW0oSWkyU+ClWu55kIajooa4cL3HSiO6c6FIFZ5cP1tAqxVKBZAR1AqeZMFJ7LmDC
IMh5x/4Cxt/NCBMl+XaClsP5DUMvlxHpsgqcTgaAuhU3w4OhwlX4uFPXuRjbDDU083r+lM9Agu9Y
0o9J/sKPlXT377zqL8yQFe5+pxfxzIfr6lGKEokkpGy/OmHZ4WNr93P484bSucUZpDkZ+5WDHfAC
tLgI9BTkeB79GeMELkq6r2vZtpjWSt6sebx8R1klEQ39oCZGjW1yKg7qRVWu1N6tIzCEsLh6bS+h
Gi4kADJr8YRk98Ed1qnNM+Wi8eT+bIpOuH8/R1wKCya49Y/l+bGs716V5SreA8xrL7HCOoj9Odk+
fb2eVRnjkUlju8ksoWW/o+zbaLN386iLLP0SO7F2kAJkfbY1tMrb5aSuWelBjrdeqMzsbiO8b/+P
bHl4JKGLyn7YujpWqvu6tLV49y8esfdJXixVBoqkJrhMaGzyldtbFg+NaFmNFmcn7blPR2rR1NR6
EdzyLZBYlnQJfA7d6DzXxprusYLP/Phfb/SSTT6AFe9zfYxzqmLku1g/L8imzgIdhY97bD0DGKTJ
k8RhvMedC3FB1GpZiJe9IgmXb3SyPbr8FxiKo9KiRP6T0PFEoEUz7UzvhQSh94bb6xSvscdg6hhU
+e9VfXcTIdZUwJHSFgO4LFiQC6oZ12TDLNUNA2rLPwriu8DznSiaUuUC1XXUQqROCcPrqCMRHTQy
7WsAbUZmMdscBlDwUHmpDOqDafH+Oi3+hnn+xRpf3Uyi3Y/BjJuiLFoelKRDp99la5p4FG/n8tor
gLtfuvo4Ul9RsoVkQ5rs4ccXGatqI6gyLbEVufpQ8OByVAVrspLdAODzWD8JOh0t/RQRT39hAywo
fRPaZGRAxvdcEvWhlJU0upuZYisjPUd/6U1to3gJdkyRQZTvpiNLs/b253RfxN2eLQklR3Z6MsEE
UAJgiu3yArEkkTMdDMKpRs+x6UHdpF3pbZidjKF57RdstCmWbVkY3jhY6gZZRKaXi3+ndbxh9Jzi
d7FTv2/SfBVKu6JF43IbSFuge+pgkWIAlNqWVPLXqk3ygxTXCMgi+hE3ULkKu+C3ZhyJGiD7fv+6
1P/DuRWFjrXA1Oe789WGskkDwD7dfoid3goq80xNeVKiawogl1NwS841EYYFZgoNYvJv5K3st0BK
it6vQPO8mwm6ILqRGA76TUCvUHl6QufpgOXFtBvJ0T15P51j+/KQBKFFf9xcHcwTNKll3Ud6XM5t
bKxRcyySV4hD5tbcgTgHZ/87g7shMHb4gW9+tHFzAVO2uTZtZ4XARbUF1+H0acFRaRQvhui1wSQT
MSmTbLlh9k0zJ0A3cWuwvkkd1ecc2Z53FnV0wJp6EU8d3GS9ZJK/b/k83VYR/G6/SWt6aayBGWqp
tv3K07C+GmeoUIvxIcfKOdWIsoRcSTodJGIGbKa9hij1LpV2eEBAX20fs/zfzfAkIN/G+KVTzJv9
4e7R38Y43sWf8neL2TqdZOO+x5n3GjrthnPgPaH9frhOJByL73QTJTKUKSmOymJtWYSuXtZcafKM
DumCzoB75W3P/GFMhoFUlAEFpbGT1fDgekTLqWkSK62Ovwi/1Q2NEkasCqhnmXRzsl8gjRKZmg5u
n9M85+bFbwPtlb37TlKs0kNN3Xa3/J/G3FEXF4kj1eJn8sDd49tR/2Gy/6XD1xJIHn6SU7izG9jB
0Zo4IE3CbZnH/crcKyUcQHsPtIM0s+bFtAxJRJ9cT0gqqThAel0KN2243vfSSKZrb+kyil3uZgV5
XQvZVMiXwabXZacoGSttRR32Yw/iQVyKJMEN6QLbZs44+7FJy69kq2ItpW47Vj8WvA+Tv0oaztJf
fZnEHJqrursuesh7IpwxIQyzM3eIXAkjkPxFTsVJMiQBXlG4ruvRra1atGPGMHyKUYZWLiUzrwr0
o5YIxG4BZTgaj1DaBJHlBjtuEJh3oadWiuQjLLIKDURNp026oWI6DjT1uKeIw3j5ZX7LCis17yPk
hBcR1KfEEK9opl7tc0ldN3ZCbeCAjKcsiLW8ygxVTkEX0LUddkuybwGUp+g1tCxofPQa7KckYYwC
qE+hg51Y2Oan/b5w1CfwQ5LNYH34TuAtZNeIETIb7tNbLXXvMeBgb6N4Cpa4EcaXSoiEqWvJUrvw
wip9kd0Iw4q0dGYH3pNruCIlEQmz8tEOTx/Pnet4dq6rAzUMwoIF9GldEbkJEJaCgKDCNHcZZPWZ
X0Q5A5IDFGAer97rQWor2UbgxRBTmMFvR4CXRASll4UpcXSk8CICMDaYc1qIHi7LdKIUqkL5dUaL
8FSqRmSAbf+KAMmxTgTdq2zHZzczwqfF169SiI/VMsd1vQvMtB/b2HFAR+wkUTKKPoRKpqlBDMo7
nozs3nVOAXu+cySHCLbgciREG3UDI3gkvK4YbewNBwAJhCDAYQFSBUW99VEGY/5FyW78maZ2O5Ox
FSHbSzwnyX6i8rD/1PvhuXrNrQqNZHG1DqudASE1vCOdckYKa50DF1PYnGe1/VfzNrm8oSEUzeHU
gPP/AvCqk9H51vq0SUzjq/uQqifo5sAIG7hQZj9y8QK+RaevvTCuSkzqzCNKvNFG+3s4W2JLS14Q
y/Dh3xangYjcYKgaZDE59WFg/TqsllIpGZRmlGnFyTRfZb9rMy8NHkBPVdvhff5fK6BXRQQkTfMO
0PAshEEa/6Xn6K4+fleTIDGhmAe9CUcYxzxBZAGPgjyZz4PcDYWa1ZQ0OXWJl86UVKZ6RFJ78aFQ
HTXl25TcMPmcJkG8PHWFjjsZSq2E3rYh2QC2C4kpZdSDTGkJvmICQg85k70CKn4FK50syltevksK
+tOW0Ik5qNQRrZOtdsY/Cuf7GLk6ULmTeRVdBF4bMKWhycG5pcmGTFsvSgZPy3FFrefJA+AxOPRO
yJdXDR9kdntnKiE/Q2mq7JP8A8nAIdYNM/xEsq2pRTHNsuzPjIyQ6VisiwPiHwVZwwMkAI32uQhC
8e0CJfKIalXSWdPYCvNOqJ5ftR9gDiIg/Av1nnvPG7PE/+3UPNgJzgr3vNFPrZNqRGEhpbPrFIv+
Jt2QF1eOghDE0zR8JpGoUT+9W4K3sV+3wgyvWPzfTQgaN3ydcWJBtfRDtZsFw3Ye5cuPVp3Y6+tD
lF5zu/H0LuFuIU1FguZaf7c14yzmb+pEL/kL0dott4mpNj4gowG7K3pb+E1njKYWudgzkpF04wA1
ZABOFZyaaQ7thFyH/exxClh0NqdiAU71K5P/J2KmHuJTAPocQmZot9Q5P0ZeSHiiOFuIuCLFPqvU
jiR6b1v/Pwd9M+z1aR6JTdpz53Pm2fwY6uMmu65TZ7sZ76dQxFLOBr5Uy13Of6j3kF8vILCryCb4
ZaU9mpNuEmhRby9W82a0aau/X+GIkRQnW7W3lBkUyzmylUnsdwJnqVOWQkH83wJyS0Dz5xytXjC/
rgFRyM1Mi2KHPw/g4AGyIHkUPrHFwih3KCc18lsAcX23uddpAV9BjMMNNT5BUNcNckwRhezvD0cv
r4/4VDOUEsr6FahCzkxbsuVHSkzOOw5NTPrLJ6R41aBaxXf/1CSv+FKiF8zlMS0sNYzzoe9XNhBP
ucV1r+bPs59HaTDSxrQrcnXrF8U1/BLBFPqOH2DH6Mlvl/AfW/2Nr0duVwrw3KRV0poDdlQ7oLz/
xaGf6OB/93IWYzuPsz/HsprmROXqz1X4qtwawBEKkBXbb3Mu4NX7uvkc79S2tlUfrsWj9O7Wa30w
uPNpV/tIz7hts9WADWJlDdpGx40vTi3cVe2Zu3C2izfwNu7HD4n06Qfb24ZRXSDR72glM92T5UMB
sJhHqXLjbqwXTME3GJAKKEwuoTGpV//kb4OgJJoiGkzVExLYKbHQrdUSzX9JKuSFlEkfgEp0VmxY
TER3iN47gPTusmFGMu8mi8tQn+ZEilCpt+j9Dvbg4pkyEHRMebOOFE4qcZJOunAAeVXXlXvDRL5a
a2j1AbZPGqhcJWZlZzkRP9WOQRjCgu4Sm3pyAB/immhp33WhpGDKiStOBPkkJ2i0+/SDaD+auLG3
KAdi33+aFkbcl/ShIreSwlOjYD0zRQXvdh2g798wVKRICwm7XUEMt8sWb59FBJkOSpWIMny2WwxG
QARGJi/a7IOazNSiGZY4ABR6J7Kr2lJ7Gf+4x7h6ErOhvB63T4DMYh/7KfDkcmpb+Ja4nXY7vUsH
2e8+m7ddM562ze7H6cqt5KFaMtIQJ+hm5uel7Ws0r+Dhvht7s37wyr769Am4sngLbK7T22pC0wYQ
f4BMwzl4H8QCte2VISsrghlvgHxc2pmT72WmICBqhrWLhJnA2Rq7JCzw03rq2qvd+ynCH7Sc6wVW
MtbeZIBvFtAD4zLo/4oirbBKec22HL+xq2GkKD4fYQtMpX4GNhe1vyHK7B6ZrsRzY20M9+aiDeD9
/islCe8RNVIwg04uv0R6kYWocEJs6inRZFybei66DE+Lza5XGmzl+Gy/QAk9PP7j0G8qvLS8WM9I
XSmYomsK3WE37K7eyt3wnQ0EEbAtu2PjmvNMu4D7EVy0dTWcU8hLQBOu5GDTmRR1MqEx+YjQPhUY
/RbzyCdGR0risnjPQgW6TeNXyd15ZQAj31qkATbM+tn48OBP5XWVccsA7oVja3sO2S0k/DjtPkUM
unfRg/E4PSruzLiBtD4tTNDBTkThyMZH23whJFXfL6vutjJD6kgo+20PXWT/4mB8K6TREj2n2q4m
E58Q9axzVapqKl0+VSUXqpZ1rYfxx+DfNEubZXYgeGRUfQb9s7ouSq81hhWh9r4PFcSHqVskEKr5
lbvoLYtLyZ5ybH0DcbUeO/5DvgRCcQ9vZ6iS5OV/4Ev8EWPTV3znkz7BsiiT8yDayPT2dkzP9W8R
++c5fbm7s0VRwhzud1UUUxlI9HttVuU8jZLLW302c7M10fT31d8BNpEujg7ItI4xjrj5/TeR60SY
++IVYjY3qHZ1Hti/B82P6isoZlPDbENVxeDVqvvpsiuqW9BFCc+9IndQgHNSyKB3u/zrEyL9i7Mv
QjXGH1YGxa/xIWeVhK+fk3x7nBUVCmOYhphimj2y+NHvbBH4+MgxVvLZnW7i+LSGwZA8VPkImJ8c
KcG/iGtXZyV8W0c7AfkVmg/ai39ipDv9fREiHcRK19sID27UHl8VCnnFg+bt7YxWpIuTfF8FwhkL
u43lWDlWeMIzXWky7DnnhDdR+yj6q5znfeKYpMcst+6MdXYL38ywnHH2M1mcnXqD0k67a1IlgMN3
7iR8gm+y7QQRqE5DqPyi/WUgyusH0yM/TP+XvABg2/OsRSw8vTeLXNoQwVIhVWbFjB42il+yc9nm
pV7l1JWRm79vW8zxfOERjSNNTuqDeIr/Dw5Nycwkmq4fs32oQzx5MvxQL00aCbhIgaDLgsRaqSGl
5WxGBWDuAB152jMiuV0plArSB6EYEJDHwxwG01lXWgbXiscvUSwWoF1T07ddIzcuRvLTn4Be/Fz+
poMn72BmZOoZr82IrSJZm3pUrWYWYQcEX/m1mrXLSIzBHNyIVkPuKTvKhpQT47GjuzfFldTGzNWn
H+L/p3h6hRasDG3VmHu4WfWm588rctlVOc9SJWSoDGcxLVmEllswlCnlsCsXETPPIehJ32KMjSQJ
vBjBGduHtJsjhKMz1K3ospS4xDMYnP5WLd1Y9I3i6TbJP3PLjwqbe+574eRyuX217zmm+YW9xfly
BJROO3dhmZZp92B+o0IpB4SXoDLJZYVqU1aX5VO1QW250pRcqKhaL4PhNR9V+OGgA1xq5RQRlVH+
K/l6Qm4oyJRdS+tmzGoQT2y+2Bfhz6EfmPZBUicjyKszJ64VvWIqGsbwTCjU/igoNwDINQE4PWUa
KCcUckNB10u4O8YrvRRWSmhCIDkOR63SsqF+akEdZqPWuLZHGV6sVMG0g/X8hXcJE2GJyo8KDfi1
woecyvbSYQYm/G5IwrGM/UsT0u/iGVOl7seBNt2Qm+E+thTrePAPYbgSl6crf7juD4IKSEMvWlrq
2WRAQw29l1Mph6vKpZQN5pDr1Hk2q4P/UBoaWvV0CSxJiPwo6Xvfw4Uap9mKKxtJ+7Eroshi7MYm
cGm1zeX/kWLLj4p1FbLSK8ZCN9+ZL/7OJoaV+x5AGlOx+pkwTGmPAOf+uK0Kec47Vk7OBENA7QPW
Uoh6HXl6EnaUBOpskOz7PpQYLbmxy3NZKPpW0wLMsiznRtZ2GdzKFQ8gmOHYvHNszYkvW6P/1xj0
rV4aKbMBgwxrumZeVy6Rgwy0z5fkeyUPaIwfqDecOjb2JRCpmy+/qba5w7Zy/PZf0rj65M2kwn0D
i+AollvX6pJkOIFXyBgRjyJjG5XKMXtLZifdxza5mla3EJEKj7Y4cf6WpVpiXu1rDRJ0i5D0mknS
/QiGvE7cJsRmeQnikbQ5m+/GIi8PxT09OeqatRwj1BkKDiaUZDImck7458bFp7dNjbPhjg+g3XFd
tvBVhUTZ1slbKpLyZ8O21tStuvcR3NNlH5zGfJuJ9KiUzlyiaNJT1+9K/hUbJVCMkXbmqGHPwcDi
urcQSQvTvi0TM3vk+2pU9gg7oDuusZE4h/GON38yMWdnjAFepOAVP/wyyZKea4RbnzDKjm52Scm/
L17oihkn//dRqRsSXDtHIP8CWrqkLifzCHOeC85f+u7KtmQFAhc7FGhvScT36ABD4/iO729k/u8k
7DwXqwMpvj7SArtdr4lpvCkgm9+pb3KkUJg654Bfbtcng37mTTkygyadej6Z/nTC79YXjdYHdoHV
3I+hB1VB6e78Z2drhxR3vWptJoizD7k4FRRYvyWMqG3CS769LYaOpaJm/pexLdPxxDQl45AdXdev
968+IbsKsqqiibtMWTqK7+zRFDnEIV5wTv8EtA2xRUx5tNMKQB4/qoXIAGtOaEnWylMdiGUHZQRQ
z2AELIQeI5ktKgzkm9RVcJHj0O5zvNqLE5cV1x0BBxw1MOJecMte5B+nwoEILwGCPb8VsQvG3n/W
k9+e6xCqWAeSkQoLmWRC1tlVAU9dmV03B64Ewwb56zzf1ch6o5R2/V2os75RLviq2P0Kscy/Z5fu
n7mB+bebdyyRnNorHP4INB7xsX23ExbYMcQ8zpJxoeH1cdCXya+1SkxzY/B47weF7l1Zlj0x+Kjs
5fQ+XJLvnmoEMlkVTIs1Bj9UJFDNdxfqai9BSvlmZaWNxCwrPOeIWA95brOwzBtp5tDgzurx5vwj
hdSG1ZwtN82d6ck2sNSjjZNcffiPPf+dbJszlkiAfll2MqRbIWZb0UVBJ4Ie5u7ymqbxwPxEfpHK
dK8ujIsK8Ll6sEYH61os+MzPATKIEYhm4mudzLWwp3pkLkG/WZFlrHJHbWbst6ou3EilDUALW+Xo
kYzo21OiYq5UgSlK2UAS6W16ZIR4Gf7YGV09AVCu0YAm/2JwMYpBy9bBOdzSOifERTnIMfCTlPhE
MqfJJwbiZafHsP5ycNRH/omvEgC4sKoTCUrJIa3G9ffr8wt48Sf1ZK5bPWCzNRjfxFzkV/qWvbZJ
FjZTF/9nA/jRJU547rdKv+rXqNJBUcetEZe9CLs9Df55htsa2psJl/kLFYnSPscBDj8I4iIU+PEB
AVgLATfFO+hk+3HSgatxugo/Os4B+T06nDS/yDnvelrD9j6uKkxgHI6baRsHbqjXRvGR93SQwW1A
toCVxhqcNDqJDtMCP/Fg+H7DwPCLlfObAnFSibh1cxrCqNPcDQUQvYStJ5GS+A6A+//ode4l16Yv
C8elyHP2q990bd2Ym5lUS3VaFIlmLB3nXXEZatCih9dUSQaSKKl59RVbx08LAAvtRQ5McoVcAOqN
NbWZiVDIEqgXMxrQ/nrtRkOsUWYbAbadQC3bSO5yIXF199jktZGia5Hcs2yObOAQ941Xo8M477p4
lkdEUZ/3K6r6R62R5gQiDefZHWeRJTLwadbacF/scsc+M9U/rhu2j8FEi1nNTcFe7uISUm4d69zY
wH+46UGPE53a/H39TbAlMWlZC9Ehld65yBtfuuJW5jtGs42bibZCYsX/+3l+L+AU3vB+fA0xZNPX
Nqf2BrADIZb/JMCcvwq9xOeieX8Vr5WMiyLwKZ20Ijnhi1njloIKL0jIHJn3krnS8X55k5naTR6w
lGfcACZ1Uq9B/5ipX90SJ8N67UK2bmXTIZAumGYQfa4gJYNhNVvaSXV+XpBI5wJc3ox3b7EdN5fQ
orrTgN6/Fd2UOF/FK9dRx6ZvNBkoqrG41W8H3OH5PbZNwrhnfx54gEpP/EjiricYYe5fuBzt9z+H
bbIZMIav9uJADO77EGTWDfRtGydbkPiXNNgPT4FGnOosj9w0SYG9X2c3jYaCalq+HTTsFliX78vZ
Vbf4etAE/Pq2NAFApsItiH3aRAcXFd2u7IOIyJHZVyoU8lpOnYVv1kFsUjdm3IRy5n63z0i7MqYn
T00iHvJFfXhIOIePftMGmZZLyxY5+fwezrDqpnsopYdewL5cARkEHlynCSluyFsrKQ8Ej6Ycm0gg
eDSLFkgDkT3Yc05UwemgxBGcqP+2fq79Z7SivDI+13+sBtOveostFOnXZwK6YQJMPjp1gR5gsHus
6Gk4AtMM+CGtSMZKjGdyYzBM2MOkovXeb7UNl7R4+N/R2kt4AKG4hJ6AoIj9W+Rj65/Q2pSSZBXL
qEqJ62XkCZIwrEqYw8uFLKmPOYbktvZyYvvkolUkLEquTjnoKRnY2Hs/YYLB2a8f7bFdj5wZGyUE
kKheVM57ClIdgQicUfDuWJnXeVEn4BeJerSp6GJqyctFtvE3X/XxkwYGsQ9kfmw+cYMh+JwHVLrb
lFA71ERFqajxSJ34oSPbBg4IsPZS3TOmHGUaWbruNxyn87u5hWO2z16JIGrmCupEmE78tRiUzM7d
ayhUOM/y04pWC/CqsFxZfP//CxZRUvan/UqG8Z05Vp9uBDz/DkAzXtdHx6bf8bqV1J2+UXDk7Oux
VnKmP61/cKrUfLEa2yBggICFDtMqYAYJgOKTXKZGP26Wc3r+JWKY3i3aqOqfWnLAPiSlCsEf5ns2
ek7Y+eMS6IgZxLmj9x99C44iJ3/VuhuTpx8voj2J6Kxyl7vf1V8FJQ2muWfRzszAgpb+LtnSHRSw
EPJoOTKy/SCcCCYnr7BZC5hU1NiIWRbX2eE76dYrlRJ0DFChrcYFeoPb+nhibOR4+YkdkKjinQ30
ETrh2GKvQKkjccwDX8uG4fRT1DvwI45uWcAo9SvB7AhjV3AhSUzgXV2cSbQtN2xN/3D4jMDeiJCP
D8xfRhdNBnv9hwpxqDcVmNVv8grMYPhC+4q0Bu2gvooMjETN3Df2JGNm+ZFeRyEVthZBZJcKRj/s
g8Pw6k/7mtFyqOG7/WkToPQ0ZdAU/OmJKjqPf9y08zN7vBpFYQ9e+bywJTszaTSixi8KiCx9Yroi
IVLchSs6b9DxEljb7Ig3GrZlq6Nts4C2a4+AzVNq3CzPWFMOtQbezt+AgIDsO5ZAOarcIzDUHoG5
GwzaCg9ZfP+dTVA4dPzAzEefAVgTjrmfSjrbN2o5HKftCc3F5y+sEcE48UPusDgGZbi3XWbcR7VP
X+e2w/Fj/THlUw5Ap1Uup/beJoFpFVvwadTPt9N23XJx0RrjLBJOUz+r/Fs/uFX5/bVPMcD/8FYh
gB0c/ybotP7u4Ql8KEdNenEcKcxDwKgCa06bsPyvHyTe7tFyRR+nC+x1WKTMIkGKIw+HEa6JemX5
EDmqzbnTMBhBQspQfdiQ+35RnFM1jBBg7YZE1CfcMrE/gNUYicyUU3E8YKxj2k7IrLcbKSNoCYVe
juZcbom6XhSzewFkHH1yNacNc/pgBLeD1Fu6z3xGOHlJCL/d0rFpcLKbcgUJn0xqq3vubNDlgAmv
zBJObsJs1mSfnscsiJf1CaTBQwHVUAEmz/czBUP/OUT4CC+uwCA55NFVmjqZejJAQDWLeAaXGeL/
dvI3Q5Y46/I+jBZq5T4jJjwjWEOVDcra2GXqTikZivnDp41obxpPL/1ZtJiiLkR5eSiT0+psiGOj
xeIgUmxewplYUiQDMdDPnTLOSrxxoLFq5CGB/ZIqQqckCxpbpHF/Pw0ketNdV7MOvsVals1coJQ/
g0ER57TqgdAqpMFOB5FzrWiLuI72I3OS224ko4YONkcuT62+gJwUBxBvmK+alPszhWUYPS7cJMih
t+0bBvyNYDdJ5lN6P8XPDT805ZN3BHu8UpBMwMb/QoruVN7PfIeK2tcWd8kpBXv3G0BY+NkA0m9k
oojyG1ZJIFfLKPWEYtwF85UrMsfB7en7mi6IZ3p6IeC8QtPXkJrnTYZp/MozWmYH/XnbXeGb5e17
dm5e3wraz+9RVBpCq7yD04Va1F0TZuMr0UkqWP8YNYRP5tCZtqWzer4KtfmHKTAHQAonKwGs86M2
v/UE+56tkhZniWfHjpKI4Bolsj+/NPnyVPAFvgOpiMNB0SVomS5J5SrIy1rKFp9jMBzMt5uY8n27
p+kS2EXJznfolw3iUBLedHU9lirtRYMEfViEwLcZHXkunV3Oh5YS/vnOBXuiDOmwHEvye0fXS2p2
+miLVDDTJnJ/7G6Hq7z2nP9d2PfLoOvrW/TZz5V0ItfS0Gm9tr5FVUG7nlj+rXD7XvrnPgx7kYta
vdBMWw3J2gQyYzhyDavDKXH6FimzaWNaWOr/oenZa2DOpPqBf3/C3j/bprf5zRM3bLSdFUpqH6Il
684tVxncVSXippalNr7Z7YCwTewDXXWt+KZUF0y4ziG/Wo12GMzB/wpeTRLJmUcBrehy/Dj4ynTv
2LSusCG/NG71EHYlT1BFk6bEtcbZS0EqL2jMD2bGz3QMjeP+cDCiNHOjT16jBqCi+mwiWzWfJcjn
W3DFKQG97U+w6x3lSwOhbdAdhnNrYV+kmTc0oIX55JZKctONb3eQjb/ew4nrTUMLHYLtxaSa37f2
yQrFJbzIrfHpDi5bWp5Ds1dHd2wxeZeXg5k++xGs7kfMevnqnGbItx766OAEwaVHmtkexWLf0ejW
co/4azrAjPu0/KUmPYl4riq2eAfu8FCpPNu4DgYi8x7P+yeJT1OY/DmZHV6+y++/IYI0ntrMdTwS
nCJsl4A3LgW2q7VLcl4/IIOhctNnf2wZ7qXdHwTHyjja83Hc11X3gnnBxIzqPBAX1AJRZnSmaOGg
7iR3C/yngplfPgpxBjbuj2WjT3F2bWVzPz8AYOjDeHuWTdy3fZVBIka8x+Ly2wMxf2Hhn0NWuGdG
r1v2MACF2PUjwv1EP72xiMSc1BdGMdEUUvSfBfhk9Qj8UcVu9cH1xS40GcPperWKpZ5tdZJ5LZE4
GYP1HujLWKOxrljsG4WwJc3mtqsYMB4KxSJskbp2ZS0uxyeBNpi3TsrUzzrOnflNnynkgB6d57G+
CEs8d0eph13rysY2lKtBy8KgOYlb4yeg7zanrJQx+hBTvm91cPr1BhIsPsYNT9kz3z5/lEGz6QRE
qqdjkcayNXSqIoYL6PX5bc/mNK1N5i6ZpO06IjAwhlI2iYju43HE2m1xtmywouhD6Wf1SG+/RJ2w
17VEqQGDNjqcL5RaW1gWduLBsm6d3Nf+0HAlJJZovLIDyPxu2nGhYF75ErnHR94st3Rj27CSpApY
zWgUAVvDruxzYXjm1tYLwNc4pApf1s47FVgn8snZ3rU/9YxOm/hN7bCDCEAeeDj4VAEd9YmYO6/M
INfN5sUvHeeWJM26ewhJ6fdfNpeaN64z2PPkW2yWMdEU+LL0ZKBCz/JTWt+znKLQAoxGLRjPgy6x
fdZ8X/aa/TlO5tEhTGsQfSZi3ePlyZcKHwadtPC4rkgSPrbaT5+5cSblVvFwuHNOUIqRlj7UQcvD
kDJ8img/iN6uS9XqFOYpfizDzzfza06s0aldgUT2OiOw1lLHXDMAVwkJE9nSi37niVjvk9nWJ45s
HEl6BOF4AdV8yy9cpVu4hJlTAm/SKdgV7sRvmwUWXnWKjUB2/+QKbXsRqUp8iscbD/G75KDcU8pd
mu8t03dkVw4lLNx/Fq3PWy1JABJREHU+m1B1EMznDF+YCHYDQstTGzm5yi3yOnjKaejvmH/ZxiIR
R4vTJzOgHiFUfnle0ECcIfUbrWHs3dakfXgnYAVC0Sb5ZXV+VPB05OjOj4M2/22Bo67Y5WCtc1/L
i70OaWSK8a4QcB85qHTtuwaxX3N6H7bdqs7FmNRwLiBJn3NIaNEX+gIRW2KSIO/ha9cTHUiTR0nQ
Q5ozLFwe1VjzuK6zGE3Pxq3pdnqpfSHbWEkQ9WA8wChzBa4HbMupyBc96TU+PCNZBANvesMC1+RP
c/RgpcwLi2T/orYp/3bdfl1SnMspoyu9C4oudCIPy0bI2z4WfHuB42Siqs3h20LelUECAm88K8qW
6iDPZxaGffhYrkHhYxh61rnejbqEMo+DJxWdHwrdhOiPb3YQli4ORmhOlIcn0OlfBfZXCVq0IFAa
QJcjCEpPuUT5RykOAvNOe0fu0yxsD5DJKAQ5pCPe/RrOTBQ8F30UmI812qHoGvs6+GkAIxdsi44h
lzdIV9/Ik4v5t6aLkfC251QVzlTlPpwbyE12vu3+MZfBEVvKwczvctjaqgWHiY5xHkzdUpK/m7FN
icanztqHHceyOyFu/55WtbTehAFGnt/fuyyEzsA9WIsJGE2CcFDDDirFITwouA3SnTGRolPY8+q8
SC9yYb1fy+9FgY9OiD3hNSP32q988CaMFmv7gUSwyPeiJJwf0V82Q/HFBiKR5VSiTfEhWfD3KrXT
TU+NY8Eptjw7sWlK+WsWFd6zq/eIRMTmUnmGU04T3GZ4nKaFVpItxkCuPPEvD9vJG+7QTeXgeMq7
NzuMayL+y7LgaEIbbc2WZDdunEwzM4X8LVpjq4RT/R/RxoQTIayoz230X756WiZEXz29knU/yjt+
JXXodZ/pgwlCEGwnIXWPQTTd86IWAYf8cW6Y8jg1Hs+ZHKOSEZNcTIm4yzrC5cm6XJihmsrQ/hyC
yuQGqYPj5SWU+O/Es2bZyswSZuK6GKsC5huvTBNaBgp1gTIUpaSOUgSYG4nyIZMdPRYhPZhwNhUl
c5M6LjbzGdt5wzGo9NNcSGKzFXvPT6+f+gBt7vAUZCX32sc1FlzTwCgU5bTioBYOf9KtzNZY6gDp
tTLPj3Fgqjxmdpm+VWK8bhKrdc6qmcVrxhqEi7aAehEt4gkLeLCi47duWBXBbwaewbqjLjDY+tee
NI9T5jMEAkM2xref+6tAYesCeBaQG9LZ9ifp99IwZAOtNmbT2GNxlozzdMEuwwsMVfWDwwUYGn38
sW9sQEflNKy2LwWFTNxkgPZI/VTo2UymD8lISd8s2vyBtryxtLD42PovCjgDhNWvodl1deJ/xhl+
JQF2OsbukjQX/hFQm+L9X6w7ApfqkK6t1501tJyip6dp2hHbBV8fL3UsLpNUrXd74hNq9U5pt9qC
pjtGjkPwI73ltOrIiPf48GkuA11lJQ6Ob7U0vyLXEJG66eYi4DNjPnTRnMJ/j7OQah7eU3SVlzTs
tjtIxzhi46FHP0o2Z8U3iMB+WbHRE11ETLGqvXQTRhWQMWYlaVeYXg8Cj03XdCrakC8lapXIwV3r
Cg28jqe5SLL0vQQhqDvCRCldtc+RhiX8vDHU+7LmbUGIJvxBCdnYrfXJJMXVQfptF3vLN/zXwbRt
FmC8RbTZQskl+FgokYNG6V2TPYrlQOHGGgBUCgO6J/vExBQxmcf4Jr87Qk0lKfs4t6K0aWd+6ee2
JrUUOCwzaVY78Nn9VUS8DoFP+yNbc2HwQOEVFlxnYXdnqRgiDAU9NBdfEpTGj6ehWfcmQnbm9Sfx
p3BZWz2irE2RAWz6E4EjYtVTXVtNVjcSFaLHm4Q8pWJ/1mLT7kIf5kfmn9Qf40wz2JvEi0rHMCAh
sjrq49j3CZmQRDBPOEdcienQi5++wtDa6JOZbCW706nAzXOpQkbLMFwRPzGRKZM/GKEXtQ3IU0SI
BYCwZaIqowSZsKYH5kRpN6m/YvqzqrhqKUKRQ4gZqUpxbzR2SxRjjYWLnix6jg1AGVXH+ozuHDnd
QCF3sqo2lLwd9u1eeGQESRFtNFCb1AFHc47B9nxKJql7uv6B/Je87tI33N5CvV6doAWjwEENhpbj
FG+BG4c4zL8tsQuAK9Pbhqg93YoSgY5YpRk+H9nD/uqm6q6Cyel5UuZvlW5RUBcqMT9u1dPn4fxG
fi/3eEnwL1Iqs9bXGTezgojhwVScu17oa0qtPuIhAzL6iBeqBQVXSO09kXkMxBgAxxMod9//PGW4
QiH8t6NOPwDYdBhQ5fHfuLLQ5Dl8/CN7PHoXPdSK7FesG35nDqbY95zwkzLulfevHgcPyqV22Wag
cUTnH7a9iHiZH8vrOTYVMqSKagCDsexKzAgtp5teAsXLU3z5y/XtO1YvjzVl5gS/z3OI6adpDNe2
2dBsTaR9HEJfkaEsix1wHCNOJcKvia0Rbli9nTH7+MKyBHhSCNpKVPUPesP+FMvFGFdbKYB3I22d
5/BtEo+5L3S0PCEpsPW/l5lqG35+vyoI7nnrVpTkjdW9M5bwP2ArA16fn1k2zj9uz4EEUiDHdhre
atdWAb+gQqytYQfRnQTc2k8/4XiEWv/cH7rgeVamyrnL9cqZG5YFgzzkDRsQFjsqtiXPmPnTtDrU
UZXpWIIKbfSTt5gyEn1N+sTEQcloKZG81GqpkpbGYbNGJmcaEOgeu1/OB8ukRgcPK+Q5gWlb6khq
v2rbB7mlUHoYbfgVseO/vdEfV2EYq+bc2ghvis49V1+Bc5v5mKoP2LP2v/3MN/n9cZwGD7hX4WiE
PbXJelDcp9NDBXSUH08UPxRRDu3gjsg+hCCc2fM6V0r3JptysGEdlpaYUeq2YfkShI6smZllTrEN
xHb2nHBZrEAjMaMxiTPAHiOdCZWrl34/WoToU3Qbd/Gd54f3C+B5iwbMadff+VU1sXqh81Eggpfc
rOSrMDiFYDHsv49FM8oFOu2726MJm3IoTy+vzgFFIf4MmPF5DalKpv6bjzoc/kYX4AxQHnLxCquY
7uZnp/FlK/0B8ewYhDNtD/XZMNWLAAZZW3QldQP3xoWkeo+l+dEApRus054SuZyFwjCSqavtEK8u
YgsMrMjeC6Q+39c1abEZs2gnF8vYwimjdkWLL0rNN52M2/XjDUcufL7UamVgNyR3TlQv/f2hOojA
udcOfOFd8Wos8+xrjRSpiRu1Wkod+AJEkH9zpBky5uRn+j/YEBKa95Wyrgf7+Q9Ml1EntqjTxJeC
xBztRJhGGsHbfMO2CL24sY2JLe08oJbO2Ietv2loHnnRcF5fkArUIny+i+rxsn4QGcZdVEdS7W3p
BBSSX7gPVhrjqAsCSev/PEKA0oeDkW002Pb2kps3mXDPdTeA755PKnw1NG8VGjq6/Bsc1EzGlvdA
nP6Qwv9HG5v5h2VlQjlkTA1PtvdC5xtvw9XVw0W62w1hxTIDKe8V8hMUG9ANRmJSL6EwRXHJG1GN
SFAA6WWSCGBOst1M1M+GS972W9lD8/oPnHirjilMKPNytto2MegYrmJ0gn6lnXU0ImpUtFytCPNb
TnmPkSzMklOkDQwrmvpvNCpwuesqnbnUn5memFicaTehsXgSnbnSupvO6W2KnWeUo5CPar6ONu9X
VuF4oXWREIKxShe0FtAU4iWpb+3ysPvrIT/Elfz23RRiduKlnvuT9a7Rx+8tuwO+gLy8DlW93D75
/6ewoHa3Ww1q5roWuLP4QKZMomiTAGvA1aMuN27jwVmLqstN6p80lJhzn79dwQyDb1A5LTePkbey
55c0l4nD/sOFdDPvsDeMCaaDAI7z824ckDpES7coPlptoL3mwIiH+6/bdlGrBOer9JwJvCxeKKxV
osW6G+fKelGdSCGv0l2XFDMqDucE0iIL/hiKhDAgc7006jhGHWqa/1/tAemtRI/L2TiXp6dRYz2T
KDFWUM5RwAtvZru+t/hv/8EVO8Eg7B+O/I0pfCM4vzqEo86njf4OYgXkl6koOH6FKaIQMoY0cyKq
rXGHbAXyY1K4iyy9iaFVtjh8+oz1x7VEM/XfbuC3+BX8QPlqcBd6vF4KWXKyFNIiimft2HIOhOuE
/uRAQEqi3VzuJEp1Q/mFu5vU4VD6JTHSQEvDZV8rEhUCX4uD3BHEY4bEkqZCceND5nfxnxi8dgpj
mmz3vLdIzj57HOplYjv6jfh0BGtw8xVWqrT3JbbUFKY5uZ4NAPrEfQ3Y8X89lWTjJYT5t2L4VeBg
NlJOeQquriXoMkt3v55Ufj2WlUIBKbY5TAQaYJxfWaQBqxWHgiVF56MywQjqF/neBqTGfVJbvUqj
VAHGXSoaw/L6ShxchCmtoV4uEwkvO+VGcPQWCmUfNAkle4tl18us/G6+UeaEKZlJcTXnBoaXrQwN
gfiXSkfaigCCo13NPnKJhRwpq7jKGtRhYDFS5l3VJdAFnZhSqviYz0NPw05FWwgzGmf3p84BLZnZ
umuU58CPIMr0W5fTZDEYUgDvQ97I/WwqspiavnocoGHfyywVhitf9mUqEZwcGRuCPS5XtAmEXyuW
U38XiuzyDSYoVIICLU5t/DDcpS0Ebi8PH1nzozkhJMClQGVsVTksbF7PXlBWwx+QpIuZrCQjKBQl
c/9xjwu4WKu1YZ66c26fD1eSTxTYqOGWF3IyvX3npgwmMMBV1uDcOAdtEO4Pqjq5HOTHWr/hib7M
XKUVEKKqGXJCDwFfWDPsABd3eNKmjcmb1MF6xgYLMOTRxatCBoI9goTGeiWPLjTCqrGTAm1/bzJm
zXWET8R9wF9rb1quUll8MAqT7UQz1UPHbFHNByZp2Rdb1KKWIEhyLwXZYJ1nfrFGijCrai1gISam
SJ2ZH6k19Uasvlk63ajjaRt17s4zbzed6B1MMjDXgrMP8F/t9Pp5gHAieZGR8nzphh/f5XYVBZiW
lPzoXPKy5JKp6CauUTdNmtiZkVitRCDVNQg9bVp+DAcBQva0iQiNbKD3C1Xph0/r6jnKuSY82t0L
hsBj5SrGXWKFMLgbAztUaT2xLqdTmKg170RfCaWA93Zoh5Fd3seNwJWLLzvHTsuHEC4Gj/2iC3E1
/0ZWmI+g0MydbIAI2oKv7pjqUhxF7xTC9Sz0cQtJ5c1IE+KjLPg8yxfCzD5w5tMGL1JJOjqSeOFh
gaMy5iwmJBgWnypLPmm8MFfQf+aq4XA7GCWmOn+MnBT+UwtakTSK/O0FS/m/lbQS53bW48wwIArb
PoPkUd9/mLsaGdMGZV4uHBO1mG4gcToJQ/DbjFtVPSJR01oc4vqz9RPVpAnT0wXlcpBQ5QHJXLSY
Rm55KEaDAhgun7CC3kzsZYlygpVbuavA3MZQa3Cyxa8p81cxAx3PlWjM6h2YhVea9/QtIYeDJLrZ
NI8JQGPbWk95jHiTZ6JHgocSESMSPCyDp+SkQ4k27DRP8jpuN5C+9YeQQZWWjnGXUbSJdYAVraP2
mONsY7hNRu0EZ2fSOK1CMaepdoUBiWJtFMZ6+UlTeu/wamDlNh6sBnrwCXScyUpiNAwBXQ3SYFXU
oKGhA9Q6dWQ84HjeacPMM2zij/671VBDrrudbTlcKRy/Ff/jzsMP25V8XjYvnBFrtTUWuKpvrV+L
NlXhhKw+V7EWFS72ih3uMrIca9ze4VgPVTP5klz3+fXGzu3A5h32G5SMTeB1VAmHvmtGL2EBVMaR
QCfOWPEmsLRs1Rdz3hXolxgoQa3uZu68vCBUme49m8uEUjt8fJECH0SXrQSesYeiBuYWVL1CnRKd
Z6eucVjnSIsZaOtRphxNIHxBW0kTAfr1WnCrOfAjIg+tBr2ndgKFSc79SHyaiYHcH5yts1+Kt0GY
bG2Bv9jAPsHF7O8cWE/WZm8WDJE3hv2/w1apbmjKHrY6rHBzHFNQp2zsr0oNP74bFHvMSmeZhveC
ziL0v/i4++gRM3OAry941DaYCKYnEvAsqf1Y0JpIPXHCsI5NY2r+bZBEn/46x0sLubwN+GGg1U2J
Tdz5oTxq0xZyZc1gFtc+bgFk17/oDdeHcMlnVAYvmiyKeTZkztJ0vSlf41HNTWBFIjynTCezxlei
BEkVxrejmNmms7rCeL+XxAdZJ/XT5KN/34vO0X/I3s5aYaQlaDdgu8lamLVT1dH1Cp7KKM+4egOy
8pxbRsO3FvSIl0VbLVrJboTcmxUBSbj8FlpEixDbLRtXsQi8VQUCgMVIN0gY0C5ur+3FLpbP3VEq
hO4Fc9QHu3bFODBcPtBHa6RqJnyw4RlT7/f3ZxyXMLaK56qy62jFDicK1B6Y53MN+cJwF6GY+Q1Y
x3vbjFBTgMyzMnk2Q63JodADXxrsTtKNjYw0se3J5PgpPzwLhu8AdisgvquZBqgJzKXza6yFXEH9
veK4mmN5wknd94H+nwJ2m9IctbFx8lCeS9bYAvNOfss4hf/GDp4HKfof9xYcHuhzbRlDcyClRUYc
R0jMFmwXUTJmTDkJc8W5TFqxDdWzdJx8f1OpM7/oJcl5qHGPVIWZz4u866C5Od6bt5WQf5t+EZq9
N699jT1JU3n5FODXYUijnWBx9HzIUyxR64hqIF4EHzuPgreM1eATZzaC6WF9CIMwYLgFxtvcTUoz
CFMnB4UMvagjsMnawq15O+NiyprN4ruCEbEt/jPYKBQot6l1pXFShaNAzpiWGuLLt7Siwn2zzoGn
gTwWmlzEFYjd728nd7F1t6u3xiFTyzfvQekpj6KlGkQajic7RmIrtDNvRtrexDBzfcRcAd7RLDkJ
PAcze69RxyV4Dh88kJ/JrCYWefYFkW9vhoXBIYQ/kPGNxwsfR3ftK9OWIhohzKyP8xermegiD6ne
2kRZph1c50Gzu7wclvI/dMnhytyoEzSfDkCuEvl90449YmTBEOMsQtLzdqvW1WHIB42nTCxGcWmB
vDgMgL+YZaxQEWcwbsxpxS124Lnyv9kW7L66HHrcDBN+hhBKfL+S9CEYQRKOcRWd9tb2vY6TGlYn
GdffxiWzQgtG5i5sdoKh4UEFKM+NEVdjX2tVqVlIsr5MtHD9xKhaRaCdvJiMDaFO8ex8+OMuvHp5
78SwPahHegs2oyqhzOWv5W3f2oE71NH+w34o+A4wArY8m4coRKTGftTcBGtWbL/hxfoIGzhnk6w2
YE9DdFvo+FSSYFYyo4fj8eAhNZWHxjgAV9zXAG7deH3xmB/LSCUNA8BLKPY+yx0Xku3T9Z0PuZ/N
ZaOC4SB4VoD4lNGcZrR0/qG9NyfACPjRMAAUn3Efl7lifxlMiSPVtBA1gEyNDujt4P1oUgvMiWje
+Dtjg1XYHR8Vfsej0u7bXK6uyfgeZvcn5A3TENQ/qaXO5446FKZv1eYA7Sq433PXuC6a5TEs7G4C
l2uIEVEbW+kNlqkQmAV00yMP15De+zeuWnaM12q7LBM0hSaImyfQ+uS1263p5Sf0N2m/67OCw0Qu
wW1KGnYqN+UhOQx0zO8t+g5ZtR7xB9kxIhiQ/B8uZOCAvpc4QUFEdX3bq9h0RRkCEFiY1iXuk2/1
ySBiX53Wsj78yMbZtxXU4kLGOdUz7SKKxJ8NDIquQ9W024sPwU9+veOqP3rBocQ7JhaUaxl8c+dH
wQnMHnJPFFOStXZf+VppgemvxF5LRbDh2z7Vc+/ZLGj0qP7RTx0tJu84EjARpPD5UKKnT8PlSH6p
UEXPCBMtTaM1irIOhpQc0m94j+7If3bcV8rcaoIlPgbXhbXzxt8e4EIDDt6Km8NJnOiy6mBli8ID
aFEjEuZHNRX1o78vqHvutFPWytkBlyZjmpjImF0deq9TAFpI7yOB+c9AeiFMWbPqUEQHI8SgTvT0
DocTlU64ddwdN7yWaFHNSg72C+VNy25V/YT9XMeSY2l1gwpJGJzbaqRuL1LqY+SUdBk8yqtDBbdi
E/9oB04xK4hLWXauFv+1YDhGOIBlvQn42DzsXFbsekq4RlapSWD4H2wWEsEnTKnkj4WogWHd0jF3
1WTBdHKoj2SX7554mo2RD+yCTwRAa8lzsRF7gv8G7OveH5Kzs6aHi0bC+iuMi5i2Pp+LLx6FECio
w7ck8bOOjbhNXR4n8BcvpiiXP2WZc1b59Quj/v+NS4ueIgoWE3GRGWk0SaHSlTO0D7D14V1JDfez
QMqHVU2igimO/HXSKM7kt9jLJK2CIOPtcKSvmD8i7sOne7laVY5F+chl85shVeKoPxi1zYtwzA5t
OwGR2M8MYnUhk3U9bsUPyoxF+/JJshM1Nih41esIUqWiIVyGyCSUAj36j98M0P6Wel/JWk2AFTGQ
DdnGIryDThO4B2CZyZAXNqzrN8oUDwjdcaoTeothuN6/FxhWPxv0ofVBNZ09xiz4RTbrxRXaCVo3
CEIpcQmgzXTr6kqSRFEEJrcY29iuUEB24b3Yi5tSbCB5hN60R63zCQ1eY4USvmJH0cOmgXpOMQBt
nDuCdssGGZMYgfZGuNCCeYcSnQKPig1udQwAM4pfUCIzUQ+WMDDDsqnOTXmaMjIurZWyfsffkIHy
DDPcZzw6jh3Hz4OdYEooLrY1YUebvPGp4L8LKvH6msH2LOAvx/dopXOm1/CBf7NgDcLgtf3WEY3X
OcOEHkEula6UbzTTbus8hEqoys2kp6LjL7dyVS1pYUVazPXjQfyRBqQCRjkiVpRkyh+hfcMnrWrC
HYyNajINTU2gvWESUTNLubi8bOH/5gEc+4ZIOGRCFzB9lw2P8lKqj9oj8nZVDpbsnfVk1YkRGSek
LeQoo45flutjbozkmbjWMk5ttUl7mqkoJ6Iea2JRONz559UmK642uqEC4W7tFGBSK/fRcWKEiLCX
goUmsl/Y0QVeMxmNavtX/j8zmAOtYtGPUUTPRl3bN5jJQp6C2f2nKSWNSDZqvwgDBxEJZmmWJuME
msRKQJdFmVnk5leIpl0mNBYxbIzbK73ifpu36dsXx8QbAtlg95tn1myNNMn2As8MLNj+4fydaZEB
zb0vTN3mPxvVV09sFR2lQqfjW4YLISmTubxBDiUHhKftJhg/HFGrqWEty/hkJ0n7buQpwMEFot63
h/x4B0nJwbfeap3NPNdznxB2Nl2/qmPWVZGMY4OvH/ZIbqTl7uU/K8X2YNoLJWlGn4LfzsQGWFh/
nz0C87Lt3uYL57/QCrcyDC2P0V06Ko8i+BXL35ZffIF1E8DLUGjsNEkWn75Y/VCLEfnPDEy2BZYJ
4hBettAqxT2Lz9n+Xn7ZF72/yB0drpvXgQaZV4voNcqwSbC+MCTHEqluUvMeieo1GQ3slO7RT4gi
7bzfHckf8Qdsdf9C0a6n3jaVhlsDSGH/V3iSU7K/kR2KTgVk99svDDCxt5PiyZs88ULDngNnVRAJ
q1zd2xWyLkKI1sIlK6apc+d6LKaiMgD526/1jvO4qi/OnSWHmgn8IA7fZo2LHlBFocPz6VUNHfnb
weWoA1qnh8yZQrbIXLbELoD3JCJ5NdQ5HtbmICdAccl4Jtdx5pUqvU3bPnn4m07Fp9RdtPQSAl26
wSeEzzsGMZxuPnGVcOagJqNQD7i0aTRffUrzoubnLyjTRlJ6pwvxt9YxSqktkVW7HW2tRayI2FFe
svZZ8zhkuJP0SAwJFfxs+Zz6tUGFMvDzXcyXIXOl1+MqlSlJtrjbye2hHPjTBUAdhEKSRUPldPSr
ZGG16XlJcIFlTGTDPVOoOsz8KIvEq/0bONIPO25hHNTFWjjMR/X3NyRM23FHEEztya1e1tDYTmXW
GtYEWVpBMxlU6G7vAU2PWhKkCZSBlFvZhsjSYZnFE2eRgB11hNNgzkAKaegX1BM1niuKXFHqNgPp
D0unKW37y8AqHHiJm2GyBgCnpEPhgBAqEZ/bcZTEbWRsIGVbz/YsxALpXhtSHRcE5oKo7vx3gGS1
remxv0MtkUtldLOAaJpqWhuv0GEQhvrKAn1tGpg7EWFGpvj3w8mymyJQAC8kIT0/i/1n6DB63wrl
FIx9SWgWG02FkMQXS5QixAXZbLkByVh2GswFzt6Y0xyGMxu0GIECdp03O5g8vEnz00w49//AtBGB
7LPVx3gxQByudY0lOyW6wkRryLUyOpVRWJHf4h1/il9oRTjcKD0mnmW/pOoQ27XU9LER16xUP5OR
mCfGKuJb2dC5Pmnj2L2J/lT/ObJWzQ9/b/TCbUcnxco7rW4mu9WuC25ev0grUp6Wa5+Q4TeQ1zj8
teaqp4kwv+lCOO5MAwICGsgjFNaulNnC9huquA8NWOqGFcLkZ5CASMLc4ghJLex8trfTYYb3b0D0
JEGotcckc8vvD3O1ekyUYTOBVIEcTjNugDHYVWI6rh/vKmC5AGPhvyxReLU5MtwQ9hAqvkmuk3Fc
IBPdCI+tQbZBjWX2+S6ErZNbukhhhTTAzms0KoGRmcQrTCuroOnjuV7on3MWJmW89P5NDBVnQHgo
REi2iu5SzgeBz/KTvsUa9mb9rE1pj+MFL0qhtKfzzra42Le0OwuffN6BZbwzHA8/yzOISGTUX5Vc
cUh3XmQZWtR1U7xaLYVeyAjBGcSKtkD2FFR+WojtNsIrXWkLJxu6reNGqwpbEqzTO8cc9DF/u0OT
y0Cnu6WA8GSQk5bgxwyMyena2KeF0oYZcBIWwn43TJ9b9p+paU0toFmlQrOVJhcSb6sBvrlMT6zS
3IqAveSC6A0IvJSpGj9LC0V1rDS16A2NE81pLkQdiTl8aopRMC5Oc3rcoBbiXry9/MftOQw3CVk/
JUu2KQM1BHCK13Bcp8E8ld4E202bJHePsk/Ki9J7HM6HYusSavtBkHmsc2+tUHETrtNz8qu9EYqU
jVqwkWus7pkw2LEhH5aK74hSIaQ72lucdK5MB/H/JpDMo04DJOP3OMJXAv+qzY4YK7BSXarE7bCx
AvreWJaMwO+oeiXDPOY9JAcD+wl8bY87LTYTSeZgxsznPEMRukf+MUHuJpEWX5hTaYB4cNyTCB0A
AWxwNcurckxOk9k5V0X8t3YdIoJkjfsEnH+Xi4bYDPuIvCAFUTWcozBX8xwKvYA69og7haualsqt
yXfebXFAJxEwsoChS3YSD5dfBatxPYIME04fqv42h0cTMtncuFyi7iOmyBS3jTNYMBg8GkH51Csn
g/azqGPiis2id1IFt9kFKuBg84L5vmo14LJJWVCz2C4w3BbvI5ngMHSjxIXu1cYjfUCmbB3u8geU
xCF8zOH4/Tc63OGLEbEZyqrWR7wKERbf8k9LgTrAbo5LLxc/aYrsNftEp2tTc47WKb5mTqscO2I9
dmy+6FQicamPVPMBhsv9Gf7iDXRDB+M2Tjt3diBlttySnwSEol88DLMUgPrJ1tuEEZ2lTM0PMeEN
aItb0YroxF8sZXkc8ljX9+hgjisgBLWmu6/k/XVpBsP2FMdk7Dt4eAYFJb7STvV9p5H56lkgnvrC
Su/rBzZXZwLpC//LEKxSSjKApOAsc8WnDNcgvfjbuAkWc4iMKsSi+c1MPkk2WDtZiZoAlI6ExCqq
fvSem0F9F0cW7GtyrxFNyb+P0EX7ykGl8YFmsJ6z1ex4GMHTdVWIPSgekF+fo+VmXNY7h6i1P9mK
QzahmYNnLNDrZyRD/CfSYk1IamaZChGg4zVKV3LneqydpRuXsZHFlbbqfZzi+qc/Av4ILjjogQfT
A8Kq/9X6WTyKnbNBez7v9nVpRMV7SutZJwhMej56aYs+F6QJmgCkJtRl5waP7mxgwoRsvP5QHQC8
Kcc7/ZdKHuE13F6/9dYLzjMH7Rk4t/prlrxZM1IXwMBODIrCqdRQfN5R7GdlRuOR5yoHggXA+Gce
U3u3ZUytpyr0wy1oRz8cJK6RryvSdK4WYzqYpvRo4VlsuA2QX9iq9ykjaN+4P+WLJoaoDUkmsxO+
I0DizYY/GM5hbdP6/KP9Dbxpi4VQS+q7aD0ksrNzH9bNB2dgzJYn2CXZc/mo6Vpq9E9mifqt15Fi
pUwOYgZfiqIQoIMnUCi7pmmfUAEs+7M/+WnL9P158hyolETZzm1t8HihGJ6l8CXe5xhlRKa/17OD
oXTVnKtImSXjJMl8fvLPPa5ADW27PXYjO7Va249sSyuM7/V8h83JGsAcupcHp8zdemVyW6audNIO
GxYu4LkQyW2On+hPX8UoxdvDuYBbTkgaoYM5j2VniPXOj7Jw3/HLlZjUbhm5bclD+68Sm/SNLaPN
AHd2Ob59of3+uQoj6Fxrfw+NtBTqIk1EgqO8DofQL/hbn36bFmM+lrUZEkB8OvdXH9j1C3kSpF9N
plpoNuAAZdNJJHprDupbuKK+EOFU2qhaTtmyawvxi0cpkFixlluFDBLic9OUAeCw7cXCzZVUN4xf
eh+ckHTZdwuXEZeH/1uRDuFOIor/TdFr9U3kWWXGIPT1jGuJgtvnHFvRww/Z0g1lb/fIh1j9wQII
HtGp/hkF8FyiSBYWU8VY70duSUoh9G6AH+s7mQqngB3kTCs7RJeN4Eqh+cAF9Lo3lObkEsS/pCBz
7Z9jNO4km/ybZYfxErwGRft+zmZ/lgfsI+3uClZQwrnYzI6+cYvGKctP/YKM+Mx95NaE6YeN7T7Q
iCO1snzsXmw/MNYFiCRSQlDqZ3CicOXzVIRUvoubIRPwDY0E9H6QClAFSQv9QxxfE4pPNbVMhPIb
6o+kAVDllNSYJBmmtXtCfSBQXAbFyWRrbe0qjNxiO9zz+6t0Ezw/mYpd67IkG520mxGSWy8ONRws
EitiUp8aw8hValJiQvWXIQVdDBvAcpXFQeTHIrAGWK4X6I1gpYLM82ZCD4poS4y/Nd8QHbgU4OaJ
9Rf8CXNSIBmfzT0wdGBTye8eXpmAnVWACDhlHgJtl5tinkGTIO3TV1RNVXVOp7DfGcCbhzffdk3+
tp4AXO2ncrm2t/2V0tZaJC9zxF7CcWCuJ1nt8jnCw0+0aIxXm6VRpJSse9Brja42CeveCNfRqcnk
AEZiDjcC1w67apAQ4UzVvGZIp5LxSjlBiQjj7pIIV69XAManmKcY+rPxKFE2bfXBxIxETzJtM/xq
3ypRsQAdDwgySqH8Ow27Of3LVsIw5hHQF1MRpiqcEE1p2k13s2Z7Ey5iH02tkheVCZ5L0ybeAa8T
36H6BxQfHfUCH3qzmkiUmPryTyOvnIYpOSen9I/8vhxNeOorssB1Il5gC/AdKuoy8js05w/7LBmE
v2WPjwmf2BMi9ItlQ9xFxnFa67kYTthCukoKuHiganOU6yxr17Ed8/dU+4/6yo6omanGtHavztWQ
jhiNJ9F8Ft1tgR2KdMv19PS+xoq0A7J9bBPLUY25qj0KaRNNdOwUSAfMybAclXfKSAuq+ITZ+Rum
EjSHm1DryW1ug2hyM6+Ym5GBxKnd4qguX6nyt8LB62c5XHOrwAGa6xVBY49H32sNicqSnV4mXXVT
h1Vev5FBlTP+eyGgGRT5LOifWsKSba/eZllgAMw3le2nDw4TGIg38ucC0CYyjnCZ+FgzcQHBZC3o
EKjFATc6todbXZQD1iUkkNnRzul+u68/EjKjKfL1OEwvMNnwphtPcHZB+OpFXmqdsp8kwzzHZdD0
vZpIC3Lfxu2KIUy1HcUarTxxlZEyhYksGJMtGVHwD6ctUn0YXeggqUKMtQVE6GkLM/mc2BhuBOuc
uRAG4eu0EZHzj0WiV350enpyKTskEpGWE8JEjioBeIwUJXv2WnqO7Z8eTDU8vXnAWiHTv9GnED0Z
2Y4p5u4hXv5G4ANtNG0J8OoTHsl4cK+sEzv9HRZP0yH4ReNqXL6e+b0AfEZthdOj1l6KtmHrZbCY
IQ2tmaAhsCpKrMW/XpH99dRzHUmYEZ2F+JIdT0opw3TAtqdD6YA8sNOmcHao1C9TAWtgltSzeYYS
mfLsh1yKQt66hiiVngUXR8Kdyy7mDjyQs3xEckpv0UFZBP4uZTNxJY1lBxkzqTO2Hl9SYsWa1emA
qwV9cRRMyITP3aXOx32cfZgbherE4jmXKGkIeQEm2h1dK+kz04PHnTln8qKH2Uom57GO2UNgyZ4o
five9E08I5X7dnhZ1QODw7+dD4b3c/+3nPOGZ0G1TxCJ09Vgt+yXJH6hL7E56ecg0FeGr6vnsloR
Pw7Ml+dpTM5vsl5BCW7D1MQwd02fkvfJP9Qte3cwMY9HuKwydLNAJhlBcPMLjlwN2lHhvy36Y0wm
tbxdgYXZme5xu6sumT2ps3gQNeZOfaXnn9RVnKnw3ZGrk4OQb4c1jcoOxbz6OTRS1v0FyPzesrKq
yJ0WPFSLOOsMKbDX3vxX/w/UIB6PdmUExtZavSz9ssj/22kFCg5EvciWBS1+qe+dnDvKi7wlVbc4
Plalma6nLdeSMC4DHZaUECs0DIi2VPECCdVhx34j7Rpuhpc+I7GOkACXXuRGpFUmEvtY9qUz9oq0
dsffV4Pl6Dmaek/QOFSfBn1bl6PN37awAEIP5BSPSifpq9pCMdCqLpHvfuoYb83eK7PuCmcfLHhP
kvvbhr1uuxwb262O21aQcpA6+BSlGy3xJ13F6hw1E8nU+1WSwMdA6pk3EO4rh91vo/iXyOHzJDrZ
1n8UbQvBvBfu39Oocktd74ec6yAjE1OTg9AY74SsqArpjDWO7EOhaVZ8gavEKwUXYtSnpu6ExpXj
pOSPpf2tjr2UhGvFlJGyaMVNWoBA8s0uO+A/UMyVG3860Og+5geVdDhQ7PCIupX6H5QH5onZKzN1
hd88s7KIYagc3Udr/kU/gdybs5Iz1EaBWCDhDf1KTwf0h3XwHusZYKV0QG2JZTtISbtwqBucFG7M
sw/OWJHkQDY3/VUOYm89xSD9PpFg3260nRCUsLlPwPzCtWB+LC1xp4pfHksRyhJrYLqckmaUmCe6
swam5DTfCdwA4LzTjY/FRSBw2Xj+zRiChi9+gEvEggeSh9Hsd+tv59B48pnPQRoIc3WyP149MeXr
YFopf/VH4VTrH8bqf4hpF5Ir7WPi1tVj4VjMzVCxy99hzwLUiZABLvXI998Cx54oOMvz0Sp6CKJr
X5oXVedW3pTuLa6aJzxttFauP+cOSDtygeGucz26Yo6erCemAO86+mTHw7UHlXsgpY2bBmezx0p+
k+o7YUxG7GoHoxc6Dw7x6pMOe5h9aum4ouvVAA5AFtPL+a4IM63Gnn/fD5dYgLxhUfcz87wS2Zs8
ckCmOJL6zkixQI4D9b0mNYu0DE2/nj5/uS4EW+ofy8ThDH/5z/WVCjcPdQ8h7Du4bolmvo8IJDJq
nzETLRLs3wmEpH5vzbZNm6WdWAUtuvMAKQNLEdxmvn9F1be8KNqDJxWx51V8rETN5RXtfpDt6uu+
TdkEeEey0dw5HFA0w9PLkC7Ydd4q6qtc2biYgV0gDwbPpvFwH4TC4gGIcNmPhkZQORdPUZaT28zf
8bLA2tZeW/atBmqvyxeksvgLtwIQsSGbUzUf9RmmmGTkmjIihFdqdmHBgj2XsOJctHzLNh4Rq2zG
6yyLfJ792dGU5t/kUxoquUP2RirMWfEAwG1w0isgBJalm1XY3UERrANbGmEIe6TL/Iz8UjzGyhTm
ySbNShjNlypoaP4a56QO/w9j4KVwnjutGJwSTVQqakybdjXLxtE5K5pVTOuSLoM0oA3VRYn+ANNc
uleCOgS4hdY/kJ9xFhiWf4vIEhycUQEik5HKxRDuZuUFu6b26xl7zkoukI5Wpwmej9QfRtu2FrDj
a5Uz1ikDYdvgqbsc3Stq4nso9FKmjp69l39c+QB/z53lEGLGCN3+st3/ghVYk6Jk88M19gmNnTqS
TxWkJGY242u4JV/4Q6O2uKJIu15X8lYQCiY2jb3j3cfQLRhkExk6IntW0Lz3+8wB9LW5gB1e2J87
r3bMqUfB6wbsJ8Y1MopYGcXSEmzKj2LYuQEJ1viyYNypoH5w64hS8aRv1Bf8n9NrGVhytuSlHZkk
F6lAtQSQ4yKJ9gDIg10J3/SdXDLjZBaFddjpgGRlBralg2ZrpZvHFiI5+pxCfxJnbP/9wmAg4D8p
adB6ZrLWANAvy9n7mz2q2olt0ex5jk3B6BCUwmITfeXeQ6ZxzGxw2MxgB2DDlvTmD0gBX2LRdR9E
z9wVKWUi1fS8ok8XeO4OtcEyETStInve0q5XIod144SyCVyx7W3A43KtXpv9acjtwjxD4Ae+uVPr
BOJqbf/M1l+5a0XP3VCHnTaOu5Qx4CdQ6Ip7vHToEzH3Rg/uAg3Ctg8TrYm6HPy6VVxTetQG3GHS
GJEkk8IAfYmdUxSXnfbX4Hr6TblvxDQCDjawOCHfwMIiJMElgv7tjJYgCVu7dp6ck9NoKQ2enXvb
vj9dwQM724+TdT1USPngOKwvhmL46IGJ3GiVAtBAArJ1pUKO79M/j9I5L0qBLG+NbVgXdtvXlJYa
UYzAbwW9y1QHFqiUjXrQkaodiUj0VOZp3FwPpV0wJ9quqqRRQSc7PAOE7FmVUNZfxBdFZmJ8vbP9
Z96XKVwQDnooZOVI/2405y30LtogloPykC8CNpTDK4Vow9sP0Pq9ctqPTSPrjMA506gRrhZoKoij
G4Cz1jDK0vhHckH2vMMGEo6elBkc+OpqnGXuWH/SfF4Aaco74OzMSXhDUZrAlkmG9iFvj0R/c8Bw
hWRwOEOISkaaM9gHw/d4iCWOzZ2cTWev2+jelaLMt5e5LsgNkBYXTAFq3ojTyTf+e/Pdnv8avd7V
YQ6bYoATZ81qqVdbsVB1V1XCfbLikU5mdDmWBys23s9Zo8hWYlyhysWi/UH3vPdr+AHVZ9wnKqF9
WI3zNb5/rZoH3+Kc74x/IFk8aAG+1FJQsGRweTm10kS6UX4CJpb2DeEKYIf+ErNgK3WlQIkaYqzB
HlLBg4ifFsiNCqoeRdXrvB4FPmui3udXjwXxuiXuuUVeZNDASUVFShvLLGjVT+ZCtTyFt6HGTHBP
b4NiEPSdCHwYwqqcWcUowzbDB/khAc9E9dtyAUcwAgcVzAcia10DhIA9EXMNPDMe4OaMvJBn+di0
t1vdLtVzPkiQ37yl0JA2KoBbgsCmzJidr66aVvz9ed1Nj0LU4SsgjOKYRgn36Yv6aERkJsMbJN8M
qmhTK234mLCY4h5cNWzNWGdlbm3OlTv3R5Q1m+2GPnQQAif2zJ9e1Qr6GXR8BTt+0Hq6lOfR2l/L
PfgCtHlrPSN3XhH5Uw83CahGbxJ4bwegIIZqc65yJ8NLFbtutwSdXGE/LfBacm/4ewzhc7xnWC2J
mcOo3b7pKffXzo7qW5l3sJR5W6aAUPrqQaCncDP+0DmNyNy6yca1FZKjU7Og1+KZXttkrSUPlt/o
MbsGKmCxsgr5/GcCYPPYqvtqwE8fQwvIdSefZUppxGzwUm0LQaN8pjvQcBf+BTbfw+LHQBGn1NaD
+ShBmZNR/5SJ9iK9a9m4zu7oO858/vTv4x8zcJVPhKQyx3s6g34GNJHVvVVoQHkE7sacEDv+aamP
JX1UkI8ce8tNPS9v+yLPK3aQc3gfYLnJXRAHMAPIChGeT412mqWuOWH2ke2eVzCTxWO7ts2TEovk
6IoRGeIWPxt4zUCnw8xjGCzXwpGm24H2X9pttoQJzNIbq+oj4HajeNt35aMoYOiimGEJ3sS8/pqm
jSC+dp0yNawdxd7b7tEbf8IX2vfSXs3DOiBGnV3gKjoGKA2RV0YQhQyfugY8maTUHzj5u0Gx42cI
ERosCRBZJwKSlFSuOFRLVlWuVRwE3tXEMFq24UnaPe6Io+0KCUKpr7OdUTykqq7qJJySG/Se5QOF
lrYxIPAE0Jr0E88hovHZj50yR8esUZZ2NIvm5zvJPgfPR5xE5kiXgIsuHSFCHtuboFk3FTXLO1u9
nuZ+nit2y0jHx697YrvuQCYeUw1aMILIBrnXz08oDO68RRpGsqurAPYBV1fYCxZVtuD/HYb7h/Bj
9jml0DKV3qWiqAQXFt1p+0gdcnmVpXwCSyUMGFNp5yCiJtOLuAAID3xfMuxUcpwYenUMJd3Y0LHR
y3pKi3OmPwPKTuG8CUwq3OB94RJ9ek+Oq/tcla2nR9s7tCr/0re3P7qSnLbWhF5T59TgHYW79ZqO
xZYwD7HwHjXKcrfAagNTId1e8Hc//00UfSj2z+1XoCrYJd7fg/xg+UzDtpHZ//xk8PCicnuMiIBb
1FUXEtxsc4+IgRUyu/IjbAiIr2eetr5WKoast2H1lOWZpnXMcyigaNrkp3nZStm0qQPXS5cMpRsG
CYMfoKdTmyg1wNt292WH6oG1/ghmRHpdRb5Btpv95yEPm+f605QUu/hYe/RZZA5+2r9LjzkfM/PU
5rg19GUSh0vujEiiWubPq9awZ4bRP2sI0nbZ/wko/Ju7gWAb8ZmZCMOzPxt2/z2sdC66TPIn0bDM
MFZ2YJzUnoBxHokR3EUV9g+zvQVyCZLtU/7CcIHuOAEsGurwto/zkKaWKaefXMGz3lWQuRnETDPw
llld0U/1n68URjkBALEHYfnizlPA8wERW0557+xUp9BiZqyKaGx+GGxgNdPbvHS0/ua73vkeUZLI
iQ4XdfsHCiFvj2AJy4rw5sTTk02mJi8BLpHOINIH6eyEKlvvDVTft2YJHapoBD2zzAFf8LKi80Ox
iVMEFNkeynQ5SZ5rTTQvJupChD2+YZA+dk/2OeU/c6QCSm0YRR3mYPBNHXxinROsB9nwMNSH/u5L
Dur4d6szUCsSm5Sib+yST096eNN1spTeKFZbxHAlbOkruVLVEBl/r8Rsy4GFb/zDs7sMNcKGsjVq
lpmbjFrTk8xwuH647w9USNjJeBhTTblo8Nr60jMO7daHjCoDrbNqaykxvULnOasKkedczH7aIsim
FkNbvc5/r7F+PrNdwyVw+Su6a/KmTUGwKoYxuz7JmL0hLNYqWkYTLTQU4Nq3zPKCp9a0KT6aWyV3
0Z33AsBEqMH03SGGtGfJ9i5UHalFAXg4JMKecd6wYlieh8QM0Oi4jyWo0PnYycjkIi0hsXyxuN6J
12zU8wEImpUK3FLnkTy0KzkyY4y+qmRtkvKNBJtuv88V+Lrnx+1kOyd0bxhL0dXKqIGibA2nImRM
CxN1GIh+tkkWrar72HwKuFh6eD0iNIq8EIbnxb/zlAANXCt3ZQigkYyHF27ZyaNpbjto0m3hTPFI
zHMpT2NCf25D/BzZaKE99o6+zA75WcxNDb5ZYgzWGUqwTvJ2ElMSWpOVoGbJrjgyj5r4usS1xZDz
/vDx1QoSS48IkY64SBk+e/u2P/UcjasEMlWifvhEGgheVVIevJ6LuknzJFrsDZIre0qlaXFX8rbF
uzlt90zbKF9SWaHDkjDuqal0fsZpva8zvRCcM8IXKeLTdLXNSObfbnukNb+YbYlwBrTgpPxy++O/
76bouz0LQ9Dvlx0iNBKeWlKcVb3HtUEcY3bVo/T112MvA3DWH8eb+qB6VqFWK+ZEDMcXhGiekkNp
Ky17ILlC79veo/UPSusMBOBU6tLqlXGQnyptGkqDeT/Yan2cnjGuVi2gapu/hOpIf7Xl+rvqvvi8
i0LMgtQZUv5Zw1k5OxIR4gUx9dbTHfDp8YSUbMl4QK++V0TKRnS5xz+HN4uT2iYPjl3j/8ocqUnr
jXvhHzvMX51mFquZg2fWzqswAWHLPkTpGDDP7Znx+Zn/ULSBTP09QPnRtyVTm6Z8nehJ6OManBBy
YNM9wEjwC+YX1+ZJHVrmp/lwJHBxdnWViTPe6rfwArVR3NHytJzLVUjWQJF1tJoaBdFBagE+pHF1
+IeC30Z7AkQ6gKQAFPeYaZCTfZ689az8oHX301i6Ca7Lq4KWjKbctC48HrdbmNu9/mgdMw6/Ezrf
NMtW/c8lATLf0uKwTFJ+DutM/epEgyySH7lxSW3Ebs+1u+jRdljL3AjtNzYJBOrpI3i7bxkZlye6
DowmAVjgUq90cypyY2ZrlOX70vLeoC/EKNsK6oawmzNVom6XtO6xodjQG+4TxL2SdHQ+pAsa4N+a
5y+t2pU4B300uGwuqDt07Kt6NOODTzwx46no4jMqY7lbjmEw2NA+caSVT8imnlskvpSzaZZ4Ft/c
zbIwSuN0xWvnmrKBe5VM/j0T6q5hVhgndPxATvK50nsnTuOw446n+nqtnKvkRnvL0cPgepkPHFAM
Kr8Z3Zo4v5ufAhVqRPpO6gjPgQqE7bnCf3AH0kL3tBHzswPgwhqtbm74P+U2o7oErA9xJEXwr2uW
a7vW0IdxR4ctc1+GHHeKP5yzncIOX3AnTGWKYCFGQ1uDgZhB5UESQy3a8fMpCgTrauz7mTozdiFD
WKYhPJhkwkWj5Ih+EiMqH48e+YU9p40Ju25exR8HdbHRWn4Fb7mXE9fm+GpjKp+wn+tcTe4L0wmj
peSzhuVWhEHCLnq7mGT+RcP1bcibmejgKDY/zjJCpbDLO3QKnG8qOG6wSB9C2DlwTuX30gPB170V
xKFjC6uRwtGSV3ifkC9H6+OLfFFtppynutb/Q2Ncwi9FkrfGdBT32P6O0ZU82BDBwpvVPG6iz9Qo
g3Icl1q9szzoU3MFUWNm/UsS0eGArjNLMvSLjioMkNkDeDQZVl6qjl3Et5XI9ne4oXrptHA1Yde/
3piesCTkwmk1gQAEewsXjCHSdJLhx2mKIQqqkUg0iNnHytFo4YRHJg8TrN6pipLTS4jHYTd73vQh
MHzOwIfUolsufbo4EJKr0lnP9o7+B3bqMKTJ2kya0xE7GnluBUTKiLKbkA3PXxj7fY+PLvoiyKbI
mbMNQc7MIsCnJM4u2XhKQ6wddsVkG7War6ScEIRmTuJfiqhYvyAy/YpZB5UpVK725UXZhBbGjcuE
bcx7PBFINgp1G3IGNMC+T8sooC10UCu48aO3eXKPai/CVQoVmf7+66x/7mmisesoMelc4CVoLTr9
Jvft7ODtv+bX4qH0jE5EOwzOgz8vKRu5gjeK/B7Bn7CXLB0960Y0ZFxGzXd0X1eoiz707SzhrF/O
LLFgMkI4/nDDlq3Kk/PR/SmmQFBM405KzkS1lSb7aHC3uyvWKdcW51HY2wLSbh0XUJwYscfHaNFn
C0fSr/oeCU3QJELosL68ySvJOIOSYIVfHJyvI5sJ3dYPGFZtrCMfLeyBygKyeGruBd9jY98KUs+g
wdNu1rVeuUEFS+v1O+pKNEhrmqCQ0XYKKCZyFhGv/bfSusmkXI+E4K95yDfXjRsTu3kHVDnJ4JuY
tBETDObG7DeQ5H4OqRQIMuUg1IZMa5uLwQ7CmRGSB6p0EeUGCaMPXEoANuVyz2EbuCmvuz2Ix7z7
g188jQ/RV9YGipVKQ3BfqSvZ4KgVlwB74daSjg6EH/OB2JNwvzpkgTXg41f08qJuCnfLDtPD1fDW
FduEnHXxTvb2c7VWdDU34U+euvFvUxfyaS4V1lo6vPLCoaJGUbqAjWnZcVp7GoTdrD6YUeP9JpjX
dus68gfmR8ppCZXS5hgIOkkw7hy+k5HS8R5bBYrusVBkzZOPZfsTkOZzKWCIQaqd9XP3UhddDYk2
Gw0mc3gZORnIVKFO94QyejFDWhRBGoGjqsOT0oxSbw6yZz7KIVDigXwag8A7PgHa3hQC84RIMGb1
UVrnL7kFptffjmGNrDlvjJIHpDpp0WkofW8RC1VpMCC08fifyoYLybCCqMjkP+fhEIz6FXTa0h7E
DJ2jC6nGBABo8c27kEk/MzfV8unsG7qBIbtrxXjpeXGJhBu6Vbbax5Isvnx6tEfih8v/NLfJAqtU
YKx0AO9sn8qMlVSmZPjYRBkNoPfZZPZCatYrP66knyIsD8A71oyfdAuKBwywPg8Q3kVZZ0fzHuPz
ChhlOqz937V2iGWo3fsQpuv5PUW7aa/C8gxhyzNqlJgXPqtTHQEv5MWTXsvDjLtgYGsNFElIYmWI
Vsx4L/Uw5R4s2T0LB7hkxJmFwcH5Rlxu6wUu34F7Bs0iMFwv2hHrgZSC8uv+wKGesxjq16nUpy+J
hbOOLC0Ft/XtOFSOAD1fhAohiHOSL+dlkaw7aOCkOuPZRPjTvywfnum9Ym1oRgGS/Au6ISkusAob
3g6t8JoHGnVSK11cWL1jYjaNx1SqgQOJ3qhb8MRCYABaOTVL2AFgsAFn6kvnN9HUj8eg6sd9OJ1x
P+K/L66EKmCR0qiwHOEbkG6FnBfaUe87zMdfx1YwmvMyBj8Ji3yXIF6RUOdW2p6KhpK6oXtgDqyi
pbeaVIKZA7IHCNEz6JINaP8tNzwIrjd40hrV96AvwzKB/EiD/yEIka33pdzS83yzy1Ls93dnODJq
wni7JuRDUyvdTpImoNFHWrbOawLek17qY9yD0xfjGp37c8Vgdx0wW5Xc0L/xiF72b0wR3L2MtjIh
3r62QgirM/eEPIo0kJvxj2P0pzfLdgRTj8b0CA1d1g2JgA49AR+Y8TfKZyRPkXq9wJVsYSvKcqkM
sYG7Oa6Uy0GIZl4ZdpYHVgL7BbjABkVOdRupBjeqk/E9grTmKyXIkUVHTJBhQzHoTm0Pu/XWUFQr
1c0T6w7Ry7qCIbQxZxfxee6gLuLBLpaiOpmZ45XxOD8OChZpFbtClCtGt1NSBuaX6CckgUsH9uZY
OeUcEjCPL92JdrQN5cboWJ4FLhoDh2b4rgsns8pCsXcw3bIVpA49D+jLMhef3eTxRaiPsOZ9Pg5w
tWeOD5QJzIhCqZiWLv9ybpLViNutASpEDgoZvr0xczmk2slshYbBQCMW3dc1GsXdgka40Dz7Ad+q
y6hkrDRC30hQDp5vpkmReT/xpM6NU6xLbUR4JjFg/0kIv6zKjLXk7yUl4e4ssJLqHYFIfwJeytg5
G+Rf0HkP/BymMFiOOIKv/LT6nlCskvBEPvn4mNkRkfLUFsyYbeAZtjpPt26pH/q/A4Tgq4SeeQ6h
nL+b6v+irlHdjdsy+nBIGYB5lumB6lxnsKDK5Q9nybtmZo+3XCGIXQiLvoS5q9ScoVQXi+xm+h44
mBnHKhUdhaMVZWj6styxRTWPbzIOLDY2S1zyspF0ASKknCFLhoiIu8/JplpeUfZ3YfVWJ6lQKcvh
BlVZ0uxlspmsV29EJrCEB1h/InRMpSdXPGP4Xv42064SZT/JWlFcvDssSJoYiB4asMDUo1jQBo88
uuvtym2u6meGmSNPt6FqCh0aRGZ7gGG/SUfrwFE99/9R9a+qMUznq5q73Vmld2Mus9733WP6A1Vf
j92mbulL8UGRnO8AnBXE2vaXfVwdY2qWORzjSMgQ75GZRkRooGRETEnDF30bXr9RGtP+RaMBT+gy
jBS5ReWlX1p0SXjdbgRtBYzxbpeNHvQOEr6DVjN+PuhTDGUsna1U3WyEsbPgHqNCP6iPU+10DgaT
6yQfKXxyISGrnKxS0Y2j8aHObbd4a758Xsz/i7yQ3ZHL6yjzA3RHleFKHd0d/UcFrvYXutt6iiFK
u3mnNTTs/xt+iEHhNkBz3Bn0zhmS5sdfHHrAcl68qKpOM59kVXPVi54bLQxQdXkrG0Oh7OxX7FDL
3L+GmigY8ZSIL4U3xl+JYIya1Gq5iR8Bkep6/YJ9Rf3kCqbF9tzxGflioTNjiNNiUh9v7ZoBmW1D
BVxTHC9RAOLHAIAnYpuqt7nf1KagoNX7s7ZyaYTaHdvBBTcbuIrVNe1k0XH1cZTB6N3CKcTKe2e7
/230HlEcqBLqOcgNUa85j+a7+Rk1l28jTA6U5FaZ0QjIsWgbuzPidoJmbogek3pTiZqGSgMK6dcX
134mWCSlv4LesNvdglPM+tRLjZSRr1LgqhslEQbCL9YlFLvFxpR6LlG3VPFkJZm9PYgNaDhLz33Z
lBQzrlLonU2zUFBs6EkCzcZXpv9lVzDAA0ZxW/dszSQefDSL24dyasax8w4xNjGFJ9ZTJIrQTOMR
TU1N508oo4GRTdRd94WBB+tV2rqlyZMVmRYIzli6Jg1qqLQRIa0XTfY6KFujg79RHBRyAaEEanO9
DXXy3Y6xvoJWBi0x9eESLcxFFm9dkFChQydGPPJMZqmYjHSem7E2ep4/yS7fvGKOIfIGja/7LFqz
5U8YTw9pETA9L6LcZYoUUAhQh4e0MQnCGEiaDfIc7RgDyVgPFxYI7uu3wdNlrC+6TgsCpU7oNLkL
JN1d9PXTNtMFr7613a8z9+wyIsu4ZGqbeI0no21WksoCczhJu8PhII+qUXP6y3SiYd1pJe2jV/9V
D1iZA0ZtAqOunvHXXxQRc+zl9Vq5b2i8AlxEUDBcW7HNLbNPGCSjAs/vspmhGYsq2M4WplwbRKbe
ao1jjSQFR2PQyr5t9eNozibIsJh4IKl3u6ODj42vPHbI75YQsJwAYIqmzU5ikpJd8EM/XW94rjSR
tuoDibLlzk4pdB6VGm2S20CIBFaBT6UefWwlLdy5MdgYWY3Yx4qhI2mkPoH8+nZksC0klWrBKXp6
3WRCuD2uSAKiixZXcmsxcwqEdAPGTjl/N05zXb/SqKw8nh5V5BsmKlCsUwMiYuyKqobnFPsUkn6j
bH9faa/QjpKYZ4b2QDX/4Sk9NIYjzWFptAMEv0PwzcBgm49iqF5pVYZFd3sqyn0ozSzOT1VI4wNQ
uqSIC2Oy8ttWN+KdV/GhlKQUKRosvEhIrDcw1TuaOkPXWi1BJ/MRWXwzVtXS2LS8oDcRBTzM/1la
0dPwX8y/HrTbWD8y/lTnes1/y2Ks/B0d+qqiTLcvC6cUm9mJi9IFIv2Zf/WE4IVEqcFaWEZXVON4
IIg0tjT7q6XPppgJijWMa7UBbl0j58n405pmFffhcOuR1yqFpbHqqWwxOXi5mPoNoAvrWzJsATfH
Uu/5QYxrlBrdLnmlg1a3s4AImwr4HtTko4czM/1g4KJqMt0UJ+HjugOiiF1M9Vp0EDYyoC1CEORD
LyadNgvHzpbtjJonnlsBUTD8Hwc3Y6LCP+VwFM5c3uEqHt1DwqCrnJuSURF05VFF3Puvh00I/SRz
sHYYAogjah7iigpoBrVi2RAuyEpS03FvRYH2AVuLuy+z4aktvFgpL4QxZ0o6nhHrYBQAUK3QDLCI
CSVYoCaNUH5WGoOlZmcsqf75ay862gyrDKYzLugh3jqkOqF90QvCCFnK/UdRg9RYmQch6X8ws8xS
UPnSWF71K0d+SgUY6BAMoPVvQfOvYDCN9oXSOW271RDWIJ0W+M441X/Ut3HRgQeWTs2JVww44PKS
f8SfISWcMvAuP13Qv5a3iKHmzmWO1jrckYWFIumg2BrB/w0w4ZbCp7Hu/4Y+Z5NrobYC8IIxc6Tx
oy40ISXeJQJ0t5kxnHCcvXO/xQOzM8ML2wp84y9v0agj12ejufvlPn6S5Njpv5aYxluW9ja3xfzE
80QSXphIDWrafqL5Y1FdbsbjkqtLaXBxIEpNbejTbPE77CUiCVYreI0VziZHOvdN+fSxpYwoCV0u
331W4c3+B9/A9QB99dytf2sdbqIXPbrtIcK6QniT1k35l3F8vmZ82JCUR25aSjBHhq6gkP5C6Z9j
LqRmi5KoR45mwMQJDXOjEd82kWW/P+68bM+xBsOTYMywiFi9XC/QFhyE2WsJvq3KrcJXYlBJQN+m
Tynj3fS9E596Htfm2qe9zcZfxTKYSwZ3ZaDY3iCBio2q8XkhwQF8Kqk2CQERys2XXWuU85+eLsui
xFloNRjd0dP6swNnRZvf2oGiEXy2Hy4feTJtA/7PfdZmNmmyYwWG1xrq4/8i4cFNcG/ht63OI+8W
pAIfTU9xqWxqNupQDdf1+s4/b13mjDSo0QyHPXWBYv2hPgi1RP5XUGF9FV0GOisV7JMlDh9yopjm
IyhsVl1jqM64O3Oc2xAr80XSb0kuu+EOO1EnBVfIsgJSGZut1k8mpXvYfMmLypreTzv+m4SYmA4o
uanweLrpLiTSyy+vfpsQ9LtLqRKDa8pTJQnFXCyVPMVWkjsMeXDLD/kM/LhOxYQJ6Kw5o8c3TIiL
+eT4JgqkKXMLaksicxgyS84TVbwr96Kfn2dgEGqpcJjXZX5XzDv1LHr2s6pFtH9259Bp24Q+BCmC
t8laVRc5MFRmsAaOF9IOulOmINsjYUxE7L8tsg4ALfoWxxxjIPbFgwpQlKzLlejnvMVrmrZicnqP
d31tTpy1d5/OxQcc79iUIqgWPwt6OpeisSDbh3PwwYw7PLpP5mxPnxFgPSbS4V0ALMCZjqv31FjA
nPmS/wBogdm+1zmU92yFweyzw7+eoTAuVx3ygZC/jFGJDx8GFyl5NcpC1mjbEw2kaxWBPohOaotb
Oisn9fkBs1JLK77JtBG1f8XWIKqNqXN/GID9ZstvtskeZUxHKwLSU/5nzzjvQs/hNoraloHCVbAH
8oLSU/eehCcYhnhad+2v9H3z19BVPmI7EnzBANkuLirBmur11wLkoV9JD3Q446Y2x2L2xzfbMA//
vupOZLqdvwqLOtl27RYF4yGpt8JRJyD+ZHFSjQR4lCgkKFfox3CeTBUWiOINYsGgRy/xTuVxK8O7
sEgio5MtpRe155RTs4JGwaskcfXHDdWq+sxVfpYITQ8OaHfsBhpxraSxLsJSvWZBfseheaweUr1H
8STgF9skDI9QN0ZpKcqEU6EQODrpeN2UJC43tu6JR7+PMMoniP7y9rYsn+w45f7ap7yioZMgg/f5
h02W/bwcs5YRUF5n4AqGfIQKgDuckNBf2XxkjBFH1SlGk+grLhm5NGFZmAFfcrAVjfN6qI99eleb
8edIAFvLIGJse344W4/qn2v1HT9Mke2xErKD/tpADXy4F0l51bhMA8WBnSMTjY+nij5ln8pVd03i
4oBF/cGAlqjmXz5Cbcanr3mDtPUxem5fKk+O+iozMF9+e7C+/MpFYUG4OuUeaO8IZCfBhE58WieU
8nMS5WH2YfxnU6AE2tBZN2k72BPTpNabtXcFOrN24VqIXn/3sQfbChIgqSIK+HdafUVz+MknPs5+
bpYV3WS8+wEe+6pExWw32J6q7bMD4u/DgtcsxwNDNOJMaWZkrjkqcR2hFjE/Cu3U0AFu8e4XjelN
iXy2BSwhbxSrC0J1mpqLkC6ds9ijp1EW+hWEdvf3ke2tjnEQLCQ780EXBhjv1Goy/uXfPHYU/IgH
pB30z2V8s5LdnF8iNRswkKDTmtKwJnSVc7AayC4P9UD0QHrdQxDNPDnbO02srEylXhrDlRPdZa6R
Wr5dwnAgSsQbnpajhZSpjq+mwWfeIawKz+ZQ37O9klMssuPqErRGD0nv5UVBTcDme6O6kIATWq+u
AZpzHYEZgN9Qdjf2EZe9aQdy0LrUZNzZyPUtKafcReeTX79iXqt8AxsvBilGsjhSTGSucM4qvxg/
abNn1A+eCtfJTtgKvFLEpBMXFBd5ARWtcU3j3eMtacLUjD4qGgVASAmSp8qxGQfju0ydMioq5VBo
/r6GDvsaf5piKBXYBDO8TxGIRRHh7BMo/0PwcRaJ2ewOCRlvcs/3XFT58b4QkKgBUNlQjwRrb1EF
RFbMEbpDZSTeSVI9ZNqcfKkgpsRg744QnnKT45wcD1mBdc9KhRehVcU55srPZ/i9W3aaqcyLq46P
bYvItartr/v5UItxYX3/t0rAv3W2mqbUsmTDF4QXl9OT//dp9wMNUJaXI1hggfYz0OmgiJE3gXKR
sk+eg/MsGnhzZL2JgG22E6yXp5vBbiGNv7EoUJD9NSNnDuq7sYdp167YMo55g38ciaQnZs3bxHwg
DD9hkuSDc5bhVddgOPRMGZWsTnzPRM4dXazybmY36z9Kfnuio8mhEPQJsWxqdXmDFnfhX9tWqyRi
hCOdBd5s279fYFw7Zi/tk1jb8FcNBpa+NekmMCcfEgWwoc9q1eXJAMtWHnLLkDnagIQ9ysZYlaaL
FI5iNc/lrw+dL4dyznhnC8e0GXzdM3SulTUNleltTt+GpzbeldNCJQ7QS9YHee4/yHRtDEzX1+L9
SYSklopFyfehV5bGz6ze1C8qYbhILSXQtAlMg94jBNq4/pJJ1auOLrVYcyahRr+l60V0ZD/lYimk
5pZly12BH+8nPuPfk6pZJPtYLoMc3ZrB75lBqPniLMj4Ze2HpdOWERMw/G9wMNmjXx6hsgJh1WiG
IKHRdbg2lK+qV5bcaTFgETqCZNsz4hAbDVp7P0569YWvIMwY5L/mXHGrjs/SSst8O5M0YvAUcQBA
2UZuWSJCm9nxTaxBOwQ8vJIUw3cQ2hPGOoWiGqzH6SZGwPimH0JHyot7upLMCVpHGeFrBywlfnV4
RpiCyZ50/+GxKoCX8IdepcZ+X1KGqeW6orx89PhGKqfwRfeTG1bqjjcYmVGagd2nFDlBqlq5B1z9
w51bJbY9kLp0KCD71Rh8nFwi/S7i+J0jjelYoKor6zx0LzHuIzzRLbQ3epP2ZYNPTGQMr3ym7p3X
cxF08W7tphF22lvzNGDM5T34dVOHyQrdOCVpZD1bIjNcurV5perRX0ISTcyfZ69X/S4ZHNSIkiIw
O0Z3XsbpDxXNE+IfIUfWCcHcQQsrat+lUUBvaj1sr9KIfzyfjZONVmpUL3o2/M3H8F5eDivpNnN1
7zA02M1FkhVc8vp9uG08rOtssZAHlp9BeImLfu0hYOUrWlZqQLg6QcPBwqUnw+D/w7LD6iJX0c69
j0bbXcrJ6cVLXNc68/fHlzI8/T+Hc2XOgD06PJLJkUrth2cnpJIfh3Tyu+ZDuenLw8tGkZ9JOcVL
UMFQPqD0lUMaFy2S8l9H65C8OTa7y3/Bml9drK42Xow+fKNsuLjzvDQP4ciI6DIigh6V9n6J2M6Z
WOtOgeZqYtBPpCBSQOA10kN2zYnxkJ7mANA1izc+gidHUWOneUuTp9V915+TeuJaXyx4fEEsynVj
1jlQymr2DZPA9CLM+8W8QjRC9o8nok9wmDq633hCYzwuydCiE6Qt+vU1s53BdOy/WRZKclUUCrXK
015YHz/hV4zSRAaJ9SLbGmKFCbgF2x0/nXJz9UlDZ7Rl4WocjvDY3KLHaX3ukzCUbxvjKtTc7QQr
UoFnucMLsE/rCYfFMd+QrjHwGca6z/DKYtxTYKZe83myDX8bp6YhJsUhvaa7dq3HHUgjwPQA36c6
qHmOugHI8MUGob3pBD2AFt3zpm48rEdCqqCvOe0U3R4NgQhX5ikSjxI5+wjr++BlzU8OwHEkscy1
iWnpdssEm0KjB0f97GJ+m5IQ1wx1MFlHCOAHwSsmNFbJMIJtd6IYXEYHcB3FCL+3mrOOdPzF3esL
HkWr0OTvlfZS8J1/qS0R7KJT0VfFGptzYhrInoCMYDTjeCrHrtHkAdEIIpox0G1ffDaxuWt8/Wyn
2a9ajBtYNAcTHi6JuyZG/hfoVNSE6/quJrCbZwEabmLPnUAhxQptmSuAqMi/VnDCK/pQ5uUt0cjX
dGCsQbmrTGJO5l5xYNkGOnSU02shRovv0Xyp0He/wj28satXaLSzbf6Do9l/Lp0Nznm02Xi0BT4C
x3MUHA+xMR4zg/nFkupPR4ji1XLdrhf/l9N1ifU4IpjnUFie+kCAljYsO1WAasMgd+12ZtsA4mFH
GZHzIrYqSR0o04sjl/SBfdMAOxUpfgUAs8IBgoQ8Y5536PfXmTfEZyqmVzyFKzzlVdTi56F0X/lt
JFOJeo4+WK/a9Qe1EwpVsu08kQ1I/pRxPs/CrnxALhvKGByDrR/Ltq2WL0ydQe0IPUBO+kPxKcRB
TvpU8D9XcVk99K6k1ZXJt5yS7avTLicm5nRpEda2DaXFxa1xWdbfQ8Ayz5M46XdCV/m9SIlsKOZ4
3SgldbxBlL+kl0EIGc7KxgocnRSxTKSK/mQEM41h7OpZcjhnMRTdK1NqxBJduIoAiIgxaqysteNF
Y4tKIU6LL+pKAT+jtlWzVtIiYsy1u4WCsfmfAcXqvcopX7vqoQGyyK7y5UtE5dnV+OJdh1c8z2rz
V7hblcssPDCqaoOf++LUaaH7pqxzQFUi9iAF00f84s0FdBdJuNeN9y1a0hkvTEafao+GAomvGtsy
2j2eA5Bk7o86JFpSWvyal188Tg+Ka9X0KfVuTFlWI3eBJJZcpwdqpF0LRQ1RnFVSdoHuuFn4UBUU
nbP04MqXLi71W1N5CW+wO1W9D/HpiVpejnd1uKrTJHG2OFzgbfdsuxybGpCXH6PWi/Hp3vo0CdYH
a9VULhbQeB9eZ7SHgCONF9j7DD2yN4E/4M1d9IkzPBj71iPCWSVsjeOvta8Ix//llLFLPIgiYcbp
HMXfZFebAsQBJxEtLlfWNwGlT0prDQCKezmTxfzmgaHovD/ItPGSsiegYuV7Xrc91Mk5+1rL7wAQ
0D8n2/RxpmQycDwkVryaQok83XcrNXWga/pOV13gTMQkP681dXu5Z8b7BjJtze2HXYgAz7yi0tgI
SW1raHvXHfONGCNP9ACHsmtvSskQMuh5XEYLhJ1xgj0XLsZodKV9Rb99GThYQquMRMu1pWQolMjw
1zbhE2aJkD+VYAqup4f8TzCcPgX3ATnKGQjwHhl9LNnjgz/8Ezr3nPYmWK1h8Pvpo5lm2gpNUuU4
Mj7G90F8/7Xj8JV5TgW3z8DTjVjzfAVcmWSmVAfXWTwK85OtMn044NwrRM7ZKHpQAObur4qrY+lE
PsWQyc3tKPiQv8JKB9YdQAFOvkCebCNI84f4hacAwWWhqtCRX70v2Q9b0ySCRzcsIz1zJ9Ubsy6C
P/3X09QURld3yVQAAlhp5L7qrM/TK06F9JL/F6K6YHaAaveBkC0daQgFAAOPpFRsSGf6PBRI1252
HmIIC0LTXr+5Z1nKHdtw+/qipWPoIk8Wzg/86pfbjcNzz6rDysg+PDLmByZYTMuDUowzwTr+e5To
G2Pp+0MJCLxEu6h1cawf8Sj9Dj1IS0c6WHEKkWHH6HNXoTtY0mqZb05Q7gm60zsy85bBvpeFW5gR
HxuVJM1LKylVB5SfEmArrvTOQRQoyOXXLkhvEsMiWFexvKBT3JseDS343OlFjoSI2O51rWU2DRLC
LCsPenFCwbIl5scTs6zuhc9RWQjrvDMJcI0008SMiHNrOajfUW4L+LNzoONfAmUoZV0eQBIMgUQV
H8Qk7hJxxJ8dXEWZNjcAFqFufDxhdeqWssce0bxnngrM+6zoMUtLEKs01VArTRzbtkrZae8PPhAB
m1lWF9dak+98UY69p5cIX0bFgw+tlMDQost/KvYvxtBmQwP/gFjAkwOj/3UIWElAFBJ2tLe9EiLP
lj6Bi0fafccZ8zsHTG51LLTLLLyidkxDLEOFF2nVIYc9pn5cg2tKjYuv6zOpDgKpBZhEnQKJv0Jg
Wl9/xq99dV1AR3AgVLKjViu8jpTjKUP3ofETQ7Oh75OFDNQ/i73Q1i8zzB4sRD81fV8M6szY3NmK
0EJf9TNBVwav9lHj3i7uUkmUl2XOnPliw/jEZho001hp7v3qVks1FVrZB/NK6KN0r8degY+BeEvr
1bswQiftjLqff4Obd46GgH6ihFxF95d/v6e/n5ejLwoskQo5RnAs08DEppYnqTfsTBwlaSaXbliI
BGa48ikV5ovzcHHv40y9iV41IPH4BD4g86eYkZ3+wrBLfa7R3b2nk2rEHwBNYMpo2E8PXrU342Iz
QyX/DFW7MZTX3A75ktH4nQNCMVNMR5UKXaT+H17nmQ5DrM7qDs2h9T/pUn+9STpHxWs0X+KlekZ0
c4IFOGWRodLhaqUbM9fvC0YhxNvZAuZJe8v6aEnZAhu5wuOV2K/raYH5MBXsy6FcX+/KxSZxR7kQ
MloOcMP8qhoXaD1YjhddPyDQ19Yr3k0rHT7XnKYofqh6ED+oWbgXSLMz/qlOTIm0sdbOiTMRcE9l
o+k+fhOxFbX/wtQ5Jes/+CWmRfWTa07dN8M3p5VQk+ShZJLBARbHnRT9/NuMu/kGNHWC07xkwqFK
Ju+FTtoyX0pr81aD6UZRzRhCieDnnFPyeriI4HAj1sY4YtaBujUmHZjpkJaPkrEd919NqKCbrL2G
SmJh8yv/c+0k0G8Qn7IgsQSxIdaQJG7lo4Dkm86LKH6dQkkskZh7/aSqNXHnPjcF1NjYXCI9JlKu
nTty1QdFYXiDQvkgd4f56HroQT6dzT08ZNO2J6p+0U4GGQ0+wrfcljdw2eeFXgeDwkNopkvfj7hR
19qs/VQG9g/O8biWbzA4590k83fatLOLqGBllDMzdJ4AsrNH7CJYGAmMDng/c6GNh1AsYSkNsQMf
XMTavss3PM/uo86ytTgN57RveZpXsIGjyIfZwBNp8q32YZmmOLSxdTajgZw/JzJ4JwXyMdtqTA3W
6a5Rv66AnJcIGBmZ/cQ/f9JWm/RukuKXYp8a4vlMeAOClJPbg8Z4ZP1HGBDxMZc7UCGZpY0N2QTr
Z73uj+6PhV42i+gLik1jqn2beG3enUqBniQaUcdeX+sSan1F3D9xwH2E/UCriyLodmjvYinuHSBr
La027dy01QrjKqgnZxzqyXMWxYsOhgAcFnvUjgy0O1TbFvkwOD59BxWuFyj1rjmr7uS4mlaJc7Tx
O4mGia0oGdRH3da5xZjn/0BYhMIZrQHzqhkVwCgvgogjB1MXx2heue24eTcohAfeTnaYCqWvpmW6
S7QrGx+2QVgQNB6vd25Jm0hvS9bagCOniJhzAFYxz/IfKswZgdCeXHMrs6fhi7zjzV2Bod17WSXF
eSE/FujHjDBuDyvF5MAsH9WheqD1Bm47GY4q58sxiFcvimcY/MZKr9HkcNNzdpC11pi9J38B2PD0
QTPOK36Fdl2o0Ww4662agBb9pjl33zaIDsigOiWirj/iUmwKvhOhEoUnU3DDi/b9swTSQpfegcdo
QianOdmJ/B7xonuW+ymza0mICn4uOaP6XxnQqIjaTD3weU0NF6Z00XSIw6wR75jL3ahS+jQ79CE1
N8w02IzDuiXmDLVge0TO97E2K8FjAnsNwIYj8/vLPy0n9CkF9dTdMF+GbB2AVCTmassVt6LiscG6
Fa2aJcmdO5zPlMMQsUB1S0WpZbVWrBb3Ax3ZryExhLpLlHtWcSOrymr7RluxdicjXvgl8wlTtJwK
7k+kTaxn610tld1JJvc3cslYviM/QSkEoQm57ZqPS8dE+UeJNOHM+PZFbr9/VQ1t4PRuhTnv5f5a
RH63Q1RYzs8MAXGjX7H9u64vXPuR8r8tbh1KiOzDBsf4QyttYY8KYjuw0OK5jhFTctnnKZiTJWxS
ffhmtyxmYgAop46tTfkNjp+plZmS+s4D9X1673pJPVOel4tjrSTBKL+EjqNb5OZEy9cPfNVKFGac
JJV691+gYtefbQ+uy6ZAAVCeWNl4ck4QWLo8NJzIBzJzIJX9Vpl4xfiic9qyqEX1ehu3WRWcS3dN
6rg7aI58fqcPOW49KE5DY+Zna56eZE2hmRHrc0Tnml1/fTCEmtdieo+T74tJj9z91g05XwmxZcer
inPq/au/drhxZgW8gC/G7zjgX6qpMH5SeOem6EApuRJJjKSeFviVvR1wCTVgTOyAEUW69eBUqw3t
NZAIE8gGYnr8GwBkOr+q0XK9g/keSGFLbHeUf9qnwr2iUOxM38IS89wv44EKNrJXIdosLtaCzZ0B
UFGHPqh4kGNmue62jBLNIM2iegffyzXljXj3/DpCiwe6ZNX6ak+rS6NB0HxUeq6aMrk1QhLjFmfn
swvjyOGTsJM9AoPtbeTDsOBKrYOzOEPOJ82L9qxGToWwGn/dk0Z7Xvp/LlarFk0Fw6WoqsbWtZSS
wR8GojV5vfhDSBzalFySjBdZ9wTEIbkHZK3G9eBTjki9Jw0eif93670Sh/FErTNdQszL+PuJthox
nsKntgjzmIAkNwgiPewUupiSN7Slwx1MfLeZZ7GryOHCXYIUSSi2DcG3JeGGF7DmqeQ5Nw0G2uGF
0tTukrYO9NSYWFWmCRAlXTiJpCsiw82ota7oW9PX28mFUrHL78Xnirvy+ALalTAWJbOr/iCtbh4h
dZm/kO8ekbdVGQ+tjd6R3WRyAJgZ7D/mcZEZ83T0VMtbksfT6JBqbF+ARno8eurC4xuBm0QTZi/6
aGMaw07UdWOy0Yg4YIV/OaB+YIHMSm/0gop3QxaB6HTLBPXy0zEypnspsqZxWjuCkvqlG5tsxm0U
Ps4L07SkAKn2t//G+7DgRF4pPDzcMKppTxaaOeyCg/MhxwgloquGrjqhgM5cKmwSJAzSDKLywgOc
hw1DTBCTGzWyepyovlHyrEZz6qLLKXCckFz4j4f+zoygDKudkxrKyu/SxY3bAJuFNvxmZFAuEm/Q
MY1Zh3Hm+aOknrJ9zEhRpuvbydcGMi0Da8WdImW+pTNvCv+HRoPRrKE3XyLUQPJqJBMYHVULv89A
aE0ZP9OPf+jVSX/Z7CQIWW+sgA2OjPuG7i0V9lU0PRRW7mj6pZ10smVJy1Sd1b8g+oPynzB9Ax2E
UNwQCklmO7jpnWeo+92PohXFjReSDuTpvchve7UD5Pw7fncp9OyNU1eCvKyDSIjpeF4ix6oImkcP
uvsDVHbLh1mTCLNVGfV5A/cCDxTyAPm2g6fsKYM1u048wA+eftqAOb+lp6jgOMNnDSiqj0KeTEHN
JwszbKUUzGJmXw31sD8HA7EwGqqme0E6khJJSMtqxU9K7DtHPaqPuFe6RZmS957YoxEjqFXsNTTP
9Z+j5sEX/E1/y+8HIPsGk0PBPyGGW4up2PPIoJLF4DZC16IjTWzKwjbylrBPtMkTNExXChT6j3NR
ANTEQvHrGSPdeSqR4ITevxlPowzHbgVZPBnvmZZqGH0L71Zcoz6yyMjxjqaBq6UcGsJatry/s7QZ
nJVKDx+MjwyKoFbdjkFxuJRL7KRsALnvgOw2CQ1HXsgAJ+36Ng9KZb067gIrrSTWqwO4ZxMsdfDx
/HbW6GUvQHcTRctNPAZnL0enuaTBDVXWMVAnyrERblXj/RX9LE19SFvLHHGuOrcIkpDM9GWEBRd2
6lnwEA3uIum+mqVZNxoCmOUg7FGqvPzMGqHpW/Gp6zWBO+k36KWALo9IqwXYCnTgYXOvxmK8gF//
RYanbB+J4pUmk/5WODnRPMaFjiamFn0geI38tCOrydZVtNcvzmTRfjiHW2rDU7z3OakrcUd124Xq
MmxiSWC8L1HqUiWnNLjdVVFxkA9IdJYLUZ0/Rfox51kOB/dYWxi6AeOHhB4CFnSjvAqlQacbxlRI
PKEJRdhPZtkHsf0Rc8nS5azZzvabFhx7a1rrsWCwBc62TebKuVOf5WdP3tMDyHpqgtMlCrPvkmcB
um8b27wm2g7zxmTOfjh5IUYfBGArHEYKg6IwoBir/m4vQVVhKoAYr2t/TQJ151B1RF9kbZV56nI5
mXLqbDB5jM2EdhG9zqcdTF+bmmYZjlkhlgdJT9lBnG9kQTcpTXhD1FOVRmyuonefYVJZhkkjgogG
gPzBTqMSMMqkjDLTPZd52uaCvuilk/kEripHKtXj0AlOoV93puWDOxdK3TKH5i6aMw8c5R07mTaF
aTcBvpEy0+Q1R/H9cPwrK4lkSHX8vUNpuzkQDhpWj8B3cvIFmyx4Q3bWWbj3rO+HL5P5uvja6q0i
WtnqRZrodgTO+oAUOe18ewWGlO/+U2agKMRGoZw45Gty1iSQ0FEFukcI/h7YulxSQ+Wy0FTMT83E
FyNYijAPp2FxYLfm7tVYqJzTgjG2YknwmU0gpP6/HxMMYR+9DOQNEebDLbkfUrcgfn1CyTGLCQL+
mUisn3enIJ0d6NaTGKkBNCEFFrFYpH5GEpUBfrDSbtkUDztjwyxvt+LFPYUDI2v6OweKfYImHs9N
GaNZQERSehIue5gFlfLWr648mcp4OnlEULPwRHi0bXRj8qlsmUK4OdjkNz30bT9/5tD3sj0rZbXd
qtuG+mgD7um28c40EBzGwSgjZE4r2artYOfJR2utpqbVI1vZjCulXrXf+lEiCdQBttO7xlGzloTn
ToSFADAfmOEVu7fdqAeDk0Z+z8aCXfANBr6rhM1NxekXe04Q1J0OzC+7z10poyXxHTZjjfuhwqwr
RUZ8t5Iq7jVG5CA1Lp6Lmh3TfXTMvp48fdStAmxj8VJQPCMnU7UPVZ2n88wO/hF9gGykn1XJnB7m
vM0FairbQ9jJZiX34N6VoAV5pzrULQLQs1vgVNiJQHnCJhUUVR4cMet0W3wPvcvPV8J1IwwzQNtr
AvhQ1TJHKgjdDbKs80jqJUzYmLNn4KREgBRtxXszhlZQNx/MGLM1Jjogw9hExvUQ5wN1SUrwclfj
LaIyjvtZFxGONHC3MMrXfx1WcDfWB/excsAPsMq3365/jaJvO2+zlITYXFUt/MNjsMoPYdr1nB7x
bHcQ/EwCcwK5uZSFqSu27L/vWEsxbYCwOLe8eVkPzduzp88l44cdS14yaMRhUfG8+Q8QlSqVmRRc
LUKV6OXvfpTf2W9XWc9lgo3nJLVmhX28XzIZ/tJa63iFo58nmA5OQdWkPEJCJGvf5uhY+CfiSZ72
qX3VwjzDRp1s5KSRTPmm2s2CnoI8l4Yw1Ew9U2a6YUG8s3GdZQa9mwQwb6lhcPYPoZKSXKSnHZPd
HA2qVL384Zw68s60waAFgVfau3C/ua030Kda9W4xdNxoeLw07iJeIAbtQ+F+2HwYaKZ0YI9mH3hK
nY8t3PsgIi4g9mOIBZ4mx0mCJLAS3IzySpwoa/Y2/ulAZWKISZ61Zo5K8uGoWUh0xXV4hYVKMOVu
uOdKYBTdTz2LrRqMgZQ8QWSQO+2nQ47NWWJ4bIZT8vasbf8exAzX/HKkTnqAHci13IjigGkUUJT4
NIfT2MiE5GRAi7Wn5x0Oa/Bfz1ADNIf27WI3B6tBQ6S6Maw7Zocw6jeBGrBpnYoybxkrM33mDOro
UV/jeNnjm3kvlwzwU0KYufy82XkBovv7JDz758SfPErTLJp6bATA4IvZcDhfgQKc/0JuMSmyQAC7
WF6AW5r/1/oi/+xhkWtUNKN/qER+RjwYZj1af7/bJYf3eXCDXgERgYaFfrW8mkb5R/06gJqJ0nsT
durwN71YIOq+PHO3t7SJK82ug8JKpz1VfxVruquhiN1zT5H4O/OOZDVh7BvGu+m6QLvhpdpAzCzH
9XtDxdNfrLJ7iM5OgfbE310uAcBjXvyhWt49SxJCzl6P9asPjMgmG0AvgiDCEyXuKJMce8o12Lgc
DPlu0aQ/rzag5CtpliYHgA/IRO6SnlWmi42w+SOKxADmlA+Egrt/VO3cgOaehQOjPF7g9VFbCHcD
uUVBMGmqHrm8gVP1GXgxWaYlGjVaLMPXljde9K9gt4IDGsEg7m8cnVcOsvbVHDmE/i3WK4XvbZLP
kgJoICBvGQy512AJlZJzdgVX3sX36bYKmvOcXpQQGRLH1ltLLsvZ0FDhf1rS5JM5qcgHLzzRt+69
UT1KAG5xCA8Qq98+72F5qucCqLTRAYOaAHUnmV27Voffgxt+TRcKNy9DaWY9+T3FU5isoY97LXhE
vaDrmPTLVSWaivLzC9MH4VQUxJeDLcUinVcLmlsnLq56Vb/QcaOxbv2Ggapo3AtXprzBqfySDrEc
PLHId/J/kiwuCGQOWUu50bekACo3QQAvlsc0/HhoKzXlNrin0hDxuDWOpdVazJla7KqrvgtF9Qxe
fNVTjKn7os/b8mpnAiFVfk8gTnHub4uXyENhSiGlTueGE2IvE9z38l/G/O5v+8IE6+oi0yIT8VxF
CiVUgMcFCavVE3CN0cEK3DajRmedjqABHKzNom2Cki+I9qRVenljfYxE2mMNyE4CqIh0shbykSYl
8sGgMmeVfbt181G4dVUIDOey/tJ1tqrnmh7VlJ/o8qMstI6Wyjavka6a+/oElWQIUn0aZSbAgQNb
cuySwpeVl969h3hwV8Nw7zlj0F7liPsHh8gJl5AUeUx1v6Y7+kQjH/sfz+KZ13PUIs0tZ78jFpXE
laleqJaUeo5z+NE1EYiGwDKRhhb1+7O9zsOdbhTT5NwMDzOgmdYJuwlGhNTXquS3Lo8fEFvWIo4K
yFTe6ZG1W3oDUUCtbGCHnUJzOpZJtnbmAP7gvV3zg4x58YuOEPTJn2bfgjM3u8OXDiCbhul5Bmf9
lvE/l9M2CD+fB7eIo7ZilLpHI3Vtc+cYFSZ17tT63/J7Wqwvg+XXTFWqVxOHUtR2bTNh6aGpNlLT
onlpi/atb6WCrR91kiEKdYHZMLRceQhfWtoB0GXiFp/Z9PUqXEAPliUdU/8b2AZ0QbejMG/OXrzi
fao7gyw0VxVnLIV2hhbqNOfvOqWlhnVQmzR9HCZ1UoApWWfqJBPXig6tssKdnNfzTT9lXeFXhw62
aYoRnkd0vT68T/UFgjfbg02xT6hiVvimQXI2EnmpzThNuNnju+xDxixErUCfLuPWAUosct/Pc/7y
Rv0epizVYwmQivC8TUD5YeNuQcGoEKvC6Khdwf50XYRmsF1ceNnaPCylj+YPp1Vx2k/EbLxGFUEV
YQ54f6BxA0+otq20pv3/tMXArqDPLpHRbjYkmnKbe9JxUx1BLooDnvMIoTI+T0GIxT6i0q4lqiC2
5KNa/h4IMxRGbnLLoHrMkXDrVglXYBwUVdbCB/ShvQmjpb0LuQWg59p8Qwb8cPqIpFXNbVFWfLu+
rq/HuzjKfMrmuYO889GBM6zPXFzI6rnO1mLBFpkaPdx7biffMd5eCfowRdg5h8Jd4nXBQaBKAuAc
lNH0SjOBhnNut9t+bmdGSYlTeFpKQxhQ+N2xsJisWhXd4xxSBFg6YleCZi9dUT8dFQUnao3TDlKc
KMrpU6ZmMaR2D+ElZAmR3xSoIC/xqNy/MBNPS0kZMAmhkhWWJj+bkkmzJ2um+yKyA1S5wjB8mK57
C7mpqoZnrm852P5fXZQScsViXwKCiNe8RBbzJ1vx3KGxdCWHgibTpkV80tdr8zudcmJlEXf5FMcX
hWCku+ufWg5AbsvPLGNhZPoYGcJas+suIY36qIONfNGVU6odF8MFy477r2VpS9TFGMYPDC+DWemU
xFfs+yyFrV+0TVj8KD8cI87xCFkqAT3p+sluTTfwoNtjMaUg8M/DVmHGoUCI8tS+WYyif92+p2pt
eG2tqwmAGSTR/Hme44iETm0botVPz4R5XEzoqkJ91usua+oRMtcK0oESpr2tgW/FYzD96zsPhY6M
B1d1NthUG4mi5Ek7pg/0yorQio0tAGH+G0v4UlGwZGjC8UmsvEJv7YaUoXcu9+9Bh86zzl745Jtw
36bggFTbhbYloODK2sWebOlnPfeFyWg6lYtLafylW6b58SXFnYEA+EqLZ9ul2CMZr1oDmLpo/het
g8qTbz3L9uSF5Cn1Bo471R5G/oX0U40aIvuQdywpertPBp6SQrjKbAg23RjambD7PvOLDDd+L8NH
CbvfRr/f2O1ABKASb0YOvv2Ad2ILFQFouDZqSGfLosoDsimbWjHbsLUUBTlKGk0T+CTacN3rBJMa
vqNFLQyLWmu1nyli/kL70MSoPkrLxs85U0mbbcidS8niUsy0KqXrQ0c5X+80RoBiCFkkJTihV996
HMQMaT/nqrLdAEF0JrBNxvZq4V0roly6GJoy7Y3Y1KFYD/CebrAOfnlUZ2SisEAsr8eC+XO8IOJ5
vkpQNCp2hudvq3nnuGx0WHuN17VvQeFNGshtoRzntTQNXPRnJmErq0dTliK0qG60KoKwewVGKRGR
8XAks15d+vI3uacAHTnq1gXjJo2tnx3mq8Ug+qLeHSbLwN27GewFyTeamAxGhMguaU3Bkm6KzQRi
3xizCUrtcG6ocmjmlUVt6eVaI2drJEFaC5fMgBpbYLhO3lA/kWmNMbCx7xIfto0Locfk1yArRiWV
DTuC+Zhny8QyEdgf9ZWeTHSC49davYExy/hrNRVI5sG3xvOnwSKxv5n09Rx+hGSZNRyXWGViQiw0
WSVn/TcmIFiA2j0bXzeM9D3Z9B+P85/7t7guZCBBbiEaHez6heUPtW5xCEp2geLD2cYZvLPuyEA3
O6zIO6aOf91gO5++Tf20nh2dc5ZtH4N32mzARWxOqvHumyvERUBNPhUU4W/PvnFcmLKepZHijwvV
2LBD9XNsikV3fAafiEy1UPvta5Dboo6VTpobLLPnAD8ZMn69KGerfTwb7qbL011wr473l3Yq+w8E
TE3ne6geNVV1149Eyl0rAc1c9mwRfBSW7ZB8/tao9joLM7s+2L6BavrlysfVkozyIxzVI8wkp71j
LXwdbzMw2CyUxkM05UGv5hZnlgt6WCoMV5YEhXKqKZpnlPCYGxHOQfFBn4lPbJ1Nqy8r0fPOt3KM
A1CalSFM7pullmolwg+FximiC9+XZu0TRL4VqhTHXbRSwwcTAYRyTs7bb3H0NJMw5ywhkOrm/yGJ
elzn8/GrdoBDApGAh2qy99kufBH3FI4s9Quap8eEHrFjXlyFzZ/577R2lUCsNw6MJ7K/XbZ56cTX
m/MISH+zjuR0pP5430+Azn+GxBZNZQ4IQbA9L/k4kih261rFuRFrp9xj4bVkuDeMsTU4N2qdVDlO
mDRWo8BVoe9EMpqEgpCJ38657oSigPe9BrEbgvrzy5mXU0qZqgBW5tzd4P+DsAqvGn5A9gCS5wep
54qEIE65KzGKAHVg4KtBnTnxnEz8CkRZ2fozfOpJPaytzJvC5mSNDZ3TTgOT5f8YTWZBEdb95ZVD
P5cmh155Aw8pc8HL6jaBF4a9bPTGlRgGc2a150z2zgGvzOxRUsnr+KfsIiph3khXYep5MGQFyLZG
PBmxKpchZMclq/OtSaglHdsnV7uNhHn/wDkyOGpaSwlafcCAz2lmp3K7o7KssXW00AXEjs/Msqqh
kI4mNfQSaxCMrGJwDKu0DA33ns3vtd8KBATYo5daPlbirrJLTTDfIKkBxB2VOks3PcE0n2u90Wbc
ltYR2lxd1dug2UOqURbQxNS8UHKzePYQfgFoztBgb6+dWfYW/12DsKeIG8orvgvd462bIm+GJbc+
Ms0fkFmSpP2S+fBgtHBh8i3COXeKsMhVMyjRAMxPPeW3oY7yiV7q/UjHLmVTyeyNoA2EKqvd++7r
T9INJI28rAPNwfa6YZ8TsoO0ImBeAlnhLHv7Oz0x38jEMLwbQe5JImlCdEwhfVRl9poQs4E3uSmK
xV6etg4xQ7aLvQgwUnjoFlw05tlkRwdMmZGBMLWPL3AsGgQM1mH0gY8X9QzUFK3p7SJVUByyQxnx
TYBoVwNU0q/8cFovjWnPogozcDhDnb/Wopt/R3f7zp/Toktcwm+esm8p1zovbSbzLuFGzd5fT4LA
gOao7jML/CVx1ohqERB5pJVGexvIYi7uru2uF9Yj43SrGdIUGRkiGGQ9hxG13Xk/O3Uy9vWOt3D8
HfKwxIoKCikbUs2geMGg1hSSgPoD+bLhi8k/vGSMmKDdWk3dHqnMaecV8LJU8H5ESr6DD9HHGn8m
q3vl6PM/iFjLsP1zG9RTud37U5ffozv6F9uCpg1Li/9CUnaNrB2aNXINDpWlosF62NOanw1+jnPq
ZqErSpdJ5jG9nxTm0v1mvA11OXE+6lNcb/vwtapRfIf1lHPGb2wQzaK3WgoUuyWSc91WRqRgskjf
O2dkA75iumiLeM/eHRhRED9XNDpdIlNJtz9Yt2Mi+oKTpiNr4iOGVcRGgZEq/eQiKZMmRmgvSoMw
eJvn76z0bFcqpVdK2eVMCVssPoxNz8V3IAbzfz1bhDkoWaXAo2fQPJRXn/cOw43IbKN0HccecQEY
1ojQbUxomyq2H4K2DS4sadkqNmN7E2dOf7lvwuK2OYNhxV/M49DYn3slKyj69gVj72WbwkAkYtRL
mTrhNONcH5xR//gY4ijk3Au97rBugd0Vz6I5glyg+MHlPrKJ6dNCz4VeWLcpzhilZWCLeBiLLRhN
1oerdc4FS7AL1An0D5azk6ORKANE8VcJaqAo+RU+xFafa9kZw554Glqs343O4x+ln6sTFEEwnuwF
/OrEuu+6h+ClgjxI6Cve+pcT5cTKT7Rqt6X847nN+CeBGrtZQ7YpQpDHkAadEDBr7gbqF+Ztyd0S
kQK2ZBvdkkpDTcXR89/msdE+c03ztgXkI8bbVM/pQwv4ei72eLqNo8nDNI0Ztbtb3hvh/ZzHNv9y
TfJdGu8ijgDHUR8Nrjb1t9fDy54Mb694KyfTIytz98GylKIQkL1U/iG2gKtuFOJMjWbJoQ7Ejlf7
NCqg+keA/1lkq6t7Gd1tyhBgJ3teiE5Gd4VqlK2k+ppULw34JKxeg2eKwmABRtPiYT9OmBt2bgja
rXBc0sW1ZHk3pUESo95tyR9MBNcqPhv7fgbMFeJI5+CSBWRHi4BoFg+anavcgwRxK8xkMjCuWKrE
c0cIgg7mwuyh5CCzK5nabBndTAJusb5Tzf4123+mMQxyvV58blMTKOO3Bg317TrsV5Cz6+POo60Z
n9aGX6SASRFB3bhYO+4rrFRSx6tJvfi6Kgmgs37dlG6/e7pyPXCEzcpK9qZ4YGnBX6DtSGxpgKhC
xgo1ccn6NbpRh4Vp5IBsO44ntuNt0eqVXmiaNqOmMnCJE+NOpVNUOioROqS2v2y9vtN4QT3LWRnO
oT+/1VhCv//O+RgIzHRmsB7ZQlv3yLQUrXH6bqjam5HJU6IS5PyRcs9vKrFeJbG/pvEMygzyiOMx
TexJdr2vWed7Kv9Pmyax0la7bHKi84HqmMhBeatIr0h7VeYM6GFa7zMDJMnMnpHVM9XTler1FP1T
kalbXiKk6/qkW8QLmn41FP4J6MpS75W7CM4t9v0Jx35L8k5/vMY0+T3iEalTR9gYhsM1LVXm/e8C
igLi7NV4oQWqdxQZJoMTsLJd2tjDHAhQ56CiF+5fsIGCbx+TsuQuS0xa8Ixn2axPtKhvXINZGmv3
yTNN9OFpoD0LJHjZKwcvG4JM6hVf3kEG+JSNYvT7E5grA5Q5E0gheJNx1vD1f2BY5Zn6VnjTb/mS
pb+w1fDcrCA4UQ71+bvxQUcYNkKpPygthI/RVhY0kGvnqQGyqhK5oDwxIn1a8iWHA1fiQ/ZCC/hM
pGNrjoUSJ8GWi2jLm29Mi0xPuZs4cGWlqt8Z+t8X0ggEaeIuoyFOk8js9ILpD1otiDRsJ+1XaoRN
nR9cN88AFm5YIVFVDF4bnk1jmPcIE/0ZBOskFj5bC03ECYKl9+smW30SjoljfR7KhF9wmlRqf8Nu
UT2cIB1Hbyh6KZiAKBMTdrtDdNbcS+kHE9jqeFzrrC2dUSTuSU4ULjgj/WvcQ7vCefPnBVRPrkoB
sLXvHsAodAh0Es1f7ZBFEo2+nJIiYXrrztUXC+rQOqYDlPwihugOoaOy19zy1wl76V5whC8us4Ck
ClOuVBgRiUbAumACJyZ/CSbI8BOMWioSfzc6sQ4kdrXffA4riR3f/T44LoUV6IwZYK55rnKv0pS8
/1tggmLRCC6PfTpg/GZPizVzeKNcpSNqQMU5DaRcU84b4fA7e/rmjthpU4CRQPgUQml1I5DFWC0j
35HRLiHYGFXTtOBxy6lnuYOR7aFwPAkce10/U4C3jg2CX9Wsy1CH7Pp3bS2TlWcBAfwHYBqCXmAq
9vJeHiRHu6WvLe//Zjz8GYsqh1M444fjgEi3MNLM5+JtSKkewcXvwKmpoumtq0nlCA5LMjpR8BGB
/2DiKnQUFgEgZX63IxNsWiy5h5Sqv6veRdhc28rFFYtpfCY4J3kBpzruufWiqEvrhM0s7nQyrgxN
CfTXR0weeRoTNCYcKLyg0/VNC0FwGSQow9+TEVzJGXbVweuAj0R9mb7binpLYhdIRhidBHsGn9Ph
5CC/6Qzdl4LZZGgD9Fp9w1ahmvqfK+02qdWXt8cMdah/057H+kR4cB05SBTE2YGXHq6H+f74FUfm
MJy+FRWjBGudjgleU4S9kqwiCAu/a1mixLpC6rwgj1N9RbRPxhyYBmNSvj+wC2RwKEEfEXscUuy7
/tOqBcEaHMikAYOq0aHoCET0rZuzg0RmqdQVO3KtM73fyTg7uO9QtERSi+sNZRZKaiXzRCNxIBAf
HQoH1InFXIiO7/IpL6HBZ3d/TdCnYr7qb3zSCM9L+afXgxSKomQpQoityU2GEIPfwJgmgY5p9j/N
zPDCU2NDmLci+2++9Ptcd4t486vC8NLtOWRVLQk51wbIuCxyn4A2AnwhKhpojUFBNlKMZpONsOlv
brHJfVMEhaX0V8TQFNCnI1QqfVd0RjqlBtPodgGDuku+QpmUOrv3ih5oTiscO+IxLN5uZWErCaSp
JUbPlL7LC5Ef0v6lGJcTGM/JFkvzW3u9hgdCJRZJSMVRon+cdmXLVikK2MhEpdY//t9U9Gc8IA5F
zTlNIlXHDXORzCHyw+ZKGZuUtPINK4MFhuJguoQK/CsmZ3tSb0J6U3AH15A5YHyRUFIdvwPZ9NTX
SAGBl1MdP8T+uFeMBuvs3up8Va0A0sEKpJKRBnOwOB3LPPNoKl9AL1iKtQEGvRW9BZMHhq2Wxhzf
+qPlmQ/HU87OjWv1bHJVx8fD7lMrh4A8/eS56u1Yd9xXS0u5nQcnhNhXS2iGlDGwnXt+1uHEVYLq
4kjp+mxbgKDMGPUDl9no7DvORlndLns2M5z5IrZMEZun9n94ORX98n66YK30uC1je7Muqn6XuUvp
/OtzNBDgHxtBjWznORDGKNhF1LRH255Gt5Edx13msEcsH5RFz7va5Av7MXwfHlc79jNCz8srav/Z
Pluz95iwxJ/jsbe935/8woH7ZIV7CvWVoLIgbikvrgVHMGfVi/nk5jxAK14LDaW3l2+pJf6fccJa
wXvHMCJVWCU7b6Zw86iRrtebINoJr9IWS+nc5wCQpKYG/LqxvDVMt9f2HdWGbMyCG26qNF6VyE0I
IKMFs6np70wHxx04Y/uLCCWIOYDd0TJr/RCWVDJ0DzLqJ6MfTMyjge5RsU4ZwQRnQHunV/HCItZo
WrHA3B/7Q8R5ZTSYGgLbc03VP4WkU4Zln1t87VU1LV3qhgBbaJGbnuCega6kPoveazO215VrLGji
vBGeZ9zhSyU5Qq5rGdx+HrBYcUEkC71VTiLBhF/vtFZwmP5sKZ5pOuylPiJoqJjiuQo5qya7tBX/
GUWu/Pp3VXtE3dnR6KOQCQ7tslYsu8kMcLjyYwbhlP8bFSraVOuIk8ZUKMakHUCjUwjmZHQnd1lv
8vwVGRGaZ9zpQiNtMrmkYfh6An6ksU2w4TC6Ffv7RJMyZp3nX3m830mwO65ymi/XqbPIbXx9YF/0
1e1lJe5LGvjmLI7ztYr0+YAwVw5gpJEeOgQmvIiJ4dwT1gz9ThGomldMp8/hvjjnk/HraJgjfNDl
J/FzE1xStLLaokkLC4Ol6HoB5WSW9lxXzNhriaTokcAKbvBFxfQIMnRIRQpONfJMpG1E8NQTkGDY
XBDd+j8+Tima1XNpSHbTP/2jKX1lhtjHkHFb7j+QHAVCMWcRhJIynEIoM3GZLdOFqClqLTtxyAKv
Y9SJXJOxvj14aVgCTwmQLUflmJ/nlKSC5LH8HaA6FpUgxwSDr5YRMkAbf/Jlmf+K+2ENkldKS0Yi
x6We88rTYjiaqp3z3D12fC8W6Q7f8pTM/fj/XKZ3AGOanrI4w1Ob3BliQM4jVkaBTVmx45W/VVi1
2l4RLANowIIpHy9ETQ6HfZt67RHF9MoFT4YUMinfxjE5S+Y6xd3GdCM+RXY6xlOItxZ+vuDfVf4C
qtrQWVFAQAZrEGwbIJc/1d0xgLcJUYPFwjw3GB+sg+HgS8+0icOKA1kyvnKR+9wMNy36Qc+0zmqv
8sXBDwSlEVMjqwuUXiYI2XKftJqMdQSzdncydZjQ6MfIa2DtrMz2fJuo/a/uEfkL/odSVmlpsxf5
kfFRvdRLJxAz49jpHTDoG+CYeF7F3jMpy7p7Tee70Cx9sfcuoiQPWzOj9YZod4pKCAb+wy6LBZPl
giaQd4vuDka7f6DvOByVHQo1ZSZ83iHoK+fWr5eLSGkfWIuhHnHZtwHO4BxsMHSIY2Z51NhQROIp
ExG/Tt8oyRc9vC5jqtaHEC/sqFHWlV5BNQ0Ig9bs+RLN5vumVvfM0y/+/XMpirucBfBsbz1ktqzX
+q97YirvQnYp0DtySYxlXpkoVREbkasaVwyhY+AC4Fbf84upR7zQxU66OZ+eH0hGE3/usQwz1Mtm
KEV1Um+DGjHIX6PafimZ/edh9vPelK9tOOHXMENKSnjrKF8HcKim2Z/zgznPXWlO9UwZ6HwyPJuh
A0SsqFLzV5ANlbACUucXjj/cmN5iA/4QuUtHmjblEf3N26IoBRgvw2cbbahrI0+tudd/zCxhH0LN
MMhvAIv7cfMqvOz2iQeJa+EhDQEXbVHaA5R70exvZ8pqHUw7KxuNFGdolhUke06nUuNZy+3OgkXD
rMbC4uz+WC5jcjqt5xAyLfBgW0J3WWsP7KiFooBE4OXin7WVrOXdjlfxZA0phLiLrBT2UTXjyLOK
jzrW5DNX8KV+Ol0ORz7uvjTo0SliPPtfVsNN2dBP30rSP1+q7p6LCIbDhqIO2O90QgMxoAfqnlcs
+cS/rOUXSkoh91Lke2hp9UHgyaPa+EgzZt3WffdHctX9uU4c2cSlm4iMaAp6EMZArxbg6oChLpCm
pbaRQPjp1xT78m+Ld713nZTVTzBYzI0BOf6sQdJeVC3Ut1mhxu1piVHXy0wQPmKSiFETJOlyfaXl
vswQl5tFN+7P6FWrjOFXmdhyAiCALJnZA2Eu0cbe85LuFD+hD2czb/AwWkChV0ELASIhJkZpVtqY
+NnWxYMCBFs6xDXKMrp66h1k6hggFVjRDnct6eZjr+yjL3UPtLKjZX63107TLJC5X82Mcgq8g/3D
cCKjUs8mUqrI3uzFQzrnM0yE57xV+lSNEruO6WTDtsu9CoeZ+vTOlZmVcZ+HarPKVnLLwOpqyUKC
FPGGqNYfCXT4Rt3LkbzOV7CqOICf5YOuwe5AdH75nPIjNhBVd9YEQtV4blJtBBetx2oN5/QX4Tjw
jNUaNInQm24NxgxesOlXRvXz9nC3J4CRqyw+VGL8oIjXvr+Gbb30TYN4CsNlFOELc4EsUtgx1mIc
fb/7ezK0hcLbsG3nC4RAc23k6ob4xn5Lo3dkUJ9mO09mz+Tb1lz+D5PJ5V7NQniXJ+bpdBV0ENND
90pILpeQa2pcubsJvRTOMjSypC6KnjRsafKHbNEi0/YhaMf+tybEEuS5j9EOWea83DckeSDd1Tg8
D3lfwQwE8y7h5BfyLA1PWWcWQmU54WK60OPAkD1NT8ifVorM0kS4t6UInITAkY2nQQnerDJ1ii7O
T5mmVpmT4pAN46fm6DgVoigH6di6IANlcZOBpDLlELZJMcgzzwj2rr8Na+PGosPoa3KpD0ab0dni
XosLhlR4y28gkVq6MHP1b+whS5x6py4i3hhSOCJCT1gxGn+QVzzmAh+hPN9hp36RGCwWgINwO2Wt
m0hkxProVnjz/rpJHGjeNGUX+7Y6P/VszqmkW+DVxwxs4jTxdX73cI78tCWeFFOyaV5+GChrxjr5
jfDy+96jsd1DV3OUzBa2Fmdr3RYfVTfgLsK0uryWFqR4N6TRorL1xNhJPT5+VlT5y6LDdbQfK8er
DYp+Oa/bgOU6bzUGWyABD0LUh1NY1j9LSvYBgINDfKUM2A0ijOJUbRHrYUXqe5ROgziNOIGXwsnT
TP0Vsqf+Z2Y9vgGYjc3y6kyNzVwy1kXzhAvWzKOg91/cReiJQoYtOuODrAyqkEcnwdP2wED58g/J
3QRrWAX6ph2H/xKLCF8WhUITutKGLXFlvwBSXTjsQiDgx4OPGL6YBdBufgpnb0blOCVSHZOp2Iz1
P/PK+32y6eG8J68f9VUvQxw6YqgsxRfp7u+AXB04RicuqOq4tu6Xev3O/SAgelkzowy/Pqmx9ZKw
Z+QT8jPMjf/QDHuLm6Jm8zuA37oYLeKJ8oAdfvwbC1Jy3/8otxS1uMSKikJYj+4dKY49ZFgs5Blg
eAyWTqWwJeM5V6m24BPBA4FGuqwqtT6xJ+XSCRVc36dJHHCnQmc4xhk+oRdh6mzc898IbBw9UDg9
POQm/XdQmqPpR1SXMjjAF4kzdc8AxUXR9r1RXJDkIh1WEDtbXza0YLZN0MsbkrQbzjuS9VShQonY
Hk84ZMdrdJKQyGCk1SRlhMUXBuKdU7PPwbNMFNfurJoMxPwWAxIpBoX7VUNwfRfVVHE+iqqbXBHK
LTbSgiU5HLc4zZgtzUINKP4Jy/n/RjNXEvEhdE7LkqhyNg0NxwI9bJfrUG6RCYuHXuJuip0kCFOX
R4hHyKWyKLCtIFK0+Z+DQLam03Gss0hNDN207pWLwjVnl/RFNQpatXYSR0BaEFN/fu95vM5fk3Sm
iON8ZKXYCkkBWzWH3suYw6ue07GKy2sTxoeVEUsOGEM3R9civYKJKPoyUJGCTruP5choQQeblxi+
njgl5uCYk2O+ebpP9IzO6J5F6GsNifFaqN74NagIywg3EBYXtCJLpyoYAAzrIAI3y6wyzZcWmVtg
lnQepgT9+fDybPVtIiVBRUvgMfwlPJuacY+8zkkvqFWUorerCgxWyeMn4z7bcwtmQSh5cQqEdL7T
H1to5lD8crR5JJiDSGTOIyB5eFmst14GNvw+Jna8ST/Sbpg9Hmvqi6Y5k1OCkbRXCYyZcRtuZAKq
43LNcvC8nohgC7vSHm/RxWeOerE1lSJv/gx31WDx4P+ST3KbN4VXzxazulpyR+EX41VM9AyN/1o5
qFfLxvFdh3+LsJLWOhKoUK3pbywmvtlrX8G7BRc2hmQYuygh9IRH41VUv8GFupC7nUM1fsSV9mCl
yLbePLX8BNMWzKpLzdm5ieUm4Gzx1e7vpEOzD6U4Yz/2lh4WSxnlXntJ90l/hiqNnv7hdIhljC4D
7FsCi+pW7NTFLTn1XfkKPUbG+rUfpcUtzcE3XzmKE7L/aCfIGWjLzvDtGRTPe3mtry6q58Ast+Oc
cmucb5vzwp914RASIOL7PD8GnilM4QiudLaM0L/HOx3sngKPzwkWdw1EXZKA2GhHWbb2EubMji0b
BEFMMl1tVjQu5wBl0H3hE2JtTldwpszhzViLvqZJEbYYt7yIg8S6WJ/dT0lERSW7gM5pen12F8V7
oaYf8UCbPs0TR29sy/ktYZZLBGwBxS688j6eX8i8oz9QW5kJ8NdQVAKN44h43W4vp19dD/IrQqNB
zjnBBAG8KTC80MAvb/XL0NFpJ161wKIUTUKTmiA+rHXgtEZZbDM18dssnnYnylNMUrTo2MqboGxP
0ZEVcTliYkP4e1TPdi8Sjhw2PzGDbePhWFFyE8nHabl9VMORik8cs6w/hBp77/ZcHdNhEwGRQhFK
3Zg2WVWt3dbcFS5ub4Cou9+PnHsxUN1F5o1Yq6yua/2jcpWGX42kRne44/qlJaOxstgkpMlksUlL
jCoql6rbEAyegaBS0UvliLeE82DDRI3wxbMtgK+1pL34bzSZMoshGwWyBn2e2LY4nfuPc8awrI3B
/tFvoLHCAt9ZK48PQ5hra4WuX18H3lphnZs+csv7GpE5ZPv3Y+bzbLLFg0uCw73z9/+Fa89ptW8h
DBLidbJaryQKLCYQJPwAnnlGy91fOLl7t5XjPVRF6XJKKv2icL8Fk8G/ND0cyOS8MWJKCpT5fS6L
/5FUP5wlaSS8zEXQXPtWieldO/rsEyhNCcFNrE1/Hb05WFqy74sWd83ZoJdi2zKwqetaUw40Pfes
ZWFPBxCVUGDZMyfaa6ovuYLezxgTq4xGB79FBqy+JqadJgP7HVKL3mbP7LHEHlG1tj0+gFxmxCNi
zLi3DBjsdU8BM1+pr0OxFi1CrARbnkjpHuTclMjIvRpEMZFfqY+Ea1P42Sh+Vj/qenlF8gxsGwpM
4VGBksuptMN/8wYQhRwINVsfGkVBvOdytk/ffX8lrGCy42NKRenTfpiLHdnootS28FH3T4/rFRrr
daZDq47Ul91zEsRYb6HU5LFqDjsP9sRpaM7ivsHKLqWrH+xyG8A7giaN3/ZIF5YuDc6evyA6k+CM
dGROMl7rwA6aGimgf6vaWjYwBAxHplWx5Gybhgl+LSYNwPTk/ll2IXoCZ6AYLu2WKbl1uICke4Lr
vhbhsCWzHn49HZv5Q+y6zs+7+gMCTrinLfgQkgLfEtyCbwfa2iLQIqSNqIMNgV4rnB8KS5Tew2Ia
TZocyLLTBk7yEqSdZggmitDOrRsJenuCPdx+8nzk0BGwEFQMK3DJcY4RpF1Y55YBBXeE5w0aDb4T
sPgO/TZc7/nTDDDahVYHF0Ejd8AReVPlTCXCIvKRu3XyxT6VuGUUjn41b9bGzVHhOvJ2uYskkPxz
8tae2Q3qA1wcNrkUAnYfKsoaSO2ZiuJ49+L+rZQmh+Vpv8x5OwvqUwWxhI4p+WGUy6gAuDoEkGuV
K+S8sp9jb9yx2E/wYlYyY8hCAEHGrSodh5UMov+DSLMA79BTCcX8ZTBGLYxdm8EaEfLrBBtusKD4
mlk8Yo0Y95L6jbKsYklfAbOFtlaT55SX31aM8BdY/Nclkef6ASGcNTJGWpJQ5BB6WsjFCYFlbVBg
lJvZaNHcJzpebEAO7O/L5RJF8K8PCNst3qyWrJTd3I1KxYi+0i0mxMHzNdFkY2j9w/Blcy0WJsaL
aV5HO09iSbD/8uxGSgi2j7GIyCF0Sas9IMN9tIO2WF9e3J01WT1yLtFHqG7uG5FmbgArxrEtjES6
g+1Y3zgNN5kTUL6yRyoTkMCjAnr11vfqV8JgzT6UZjAuw3kgiPXPaWkYSZgRhQ4cHk5NayNfQmcM
RW+HPw5SxhpCW34YYxX+LS5KynyYQBjzKe7c7brt/REx7cCo1I3bHSkHf/tJojS7iXCkV8mEvmi7
4SmTl2h5RqvRYTHlRAFapy8Q3cJr655gvowYhBEKbFiaReB9EmfxaIZqq2vWjbmFSJLS+Zcm4NY8
0hIkO74PUd9LA+tEU3v/aesk9QeVL8Igpw/sYNiNG2B3KdhyRd8YToAKjzEPIkeT1/UI+2SVS6nm
ctTgjT/pvl3JEAD2P6zRtcjtmX9ayTFLMys98KJ6GE+8A6buSnzs3sMJRFuJrRkVtaKMXlwyTXWj
xm1P31S4v31Br0fKVmum/2+kN4pu3ipTVXVKAmsHriaYi/KHeFYerwtRXXVLH2hPskrm4vEfTjm6
uf5yNhWcrNyiNYSjE9yEPUe78zeLj9JbkrgKaKadKpeQK5+7ZiTtj4DLf4qQM9snqXJzvReKrHqI
jE6vDw73owQBoFm8/hci+wrN3FYdwpu1vZ+2gVUdcFpI50CmBY70RIW1qx/7tK0q0A/yttM2HMI8
Br9MvepSUaLSEcy0MCu6n5RS24E1BYp2dXH82Ncr04a5imA9VfHd8+zYYUgorArDMLl5rqpYjbJy
eJTpOhh+VbZnIt0KbfhsCo+Arl1dYmORJ/VJbd1XnrMIeaPirhiS7O0N3vbb7aIlUshrPC6lg710
JMkdHOwgOrIdbkAtZNEkPZieTuEDTNkSDjyfIw1XYBA+uYXvG/dtHtWZQYRMj6BCKXR07ew6zyXU
68aHHA42O07kPFyaBnefD/IAVzt3DdjFPpssjxiYsmfCtKQi6LjPyc0cbDZ/9pUEJ9w7o8HYhFZ4
gdQ2QHi9BFE+BDXHnIw0rbqHrORH7aM5DumG+4cbp5wD197I9sqjHPeGYgN8P0i2JiCozSk+qwHb
MhPQxAWlRQU+rkE268xut4vbIXqQ4HcokDcb9r/aJeKdA+Jp9Lulh0c1YJiVSSJLkuPLlvcBT8Tk
S6899XfqmaM17+hXdSfFX+SlUo5GVO50o+yUH5qVdnUDf/82NWoYddxxzPkcdK86+qhW9fuBvvjZ
q+cSrbNxz5NGfNwa9iPFImPtUIS0j4mgWFBlH7+FFr1kec1LQP0xPpdz8hhhMbdsq8BUySf261b0
RlVZLYgzE3AzV78R5OsuIyzvJoYloTPMC3eS+nVx9s/L/ULZJFnxzEshmamgrpBWKlUqwvcJwyXV
lhQeoYdvCrXCYiGkT9SCFTCVNlUryWmB96hcyX/EExKqsBVFRp5onQnvSdDp2eRSMvdAKhYT4qT1
eTcERcu+WxhWhnV6fNgASdhe7J9g0919KcHGKCEtVANpyoEAcEnTvFG2MZMajqCisP2bkv1P1zEh
3WdITmX4cjhCc+Hw0hqoWP+IF+fIWIY7Rdistek3269LsF+Mz8g+oMWrBIGiPuYHhR88e+SDJkBI
Nod7pF6zqALCUqx7OrNW7ReUUDZdT6a6qCrETog/BTW6Nn7xY81Aju0/Cq/vAXarbIzuGAf6kz2G
PygaMEyutv8GkNKPMNUzh7eI8A9NDt8wRR+ZmTBaIzDwsHLR/6xkGuqLhN26zrM8dX5IlQ163OA0
rop1Y1fWWpWqqxynooVcoq32N1B20iPKAAGCxn/7VbGK88xIdcVw9UILhYxDiJMB7OaKTybH8aNg
AYPTvh9YjUVyQ0ERMwl+YwWiMPZHOWre5gzsm5bMb6OdFnG4Dmqf9R9TLmp6tEUoSh6SoQAgyGED
lwqspFP81OJQ3SNQz7q2PSkA00wT7FuPbs+cB94XpjvWyhGJcffGvwstS56DVW2OqsnISNB7sy8p
LLl/++kwMGLURSfukGrTdlO/VID5IwF1vQQ2sgoZ9NlYiaB2p9hETfpTDino4fB+ERrrhCD4c3Nh
WknqM/NLXQf8HdZIr1G4a0ajVCu6nbTDjhujS8sB14VZC8NGsijfTgIXDdu4DH1yvw07fNHJ9TgL
nIqYXwTe2iJt4TkebamR79MpNXQPMAMUxOx9qqippsDPPuO7t5kVio3NOWUT9B56QF+7HDTI0wMb
nFbsudBIVW/78+zS4/KMnLH+w8ignycB2F1jABIds6ZUvnGGLLy7ehMCVp8nZhLsn4q3QqNeHqxm
lOD//y1Iy5Vv93QEUG+p0xukIgDItFxoi013FyJH8dQ5Cx++S3Zl54dtN1ffD9t5xKcQXgcMmSXX
9SU8IkgEhFyojobfoWV9Cx+jnWNQpGgJL91MFXZlzFnbd+CKZiOumolP4AavbWoGKpf7RjZQA83g
m4ZT/nLUzXngyAg92zXV90oLQgJ6nfFcMTX21Ht7axI700N0ORK+SlCKg4H6ZUWjXdp2X6wvSxiz
Zv5fZVEC6hllFkw5RMXcetfUibr2zjR2og4GhH64jRXY5VCh3cuWUO6IsADtlbiWyAETtm0+aPgo
VKGP9AWZ6c9ArxXKuy9LnEpaXf9UKKjpDGfVC2FXDGCP9gmhllyGt5BurNNZlodK00cNECX2Go+e
QbGFKbrI5oo2RZ0/FfqSwGPMFhQn1WsrKxGpFRD6qsG/Ep3+039Q7M9Rq6dFnKFCthN5fQLY9qhu
FE/iGVZyywZnVsJKgFKHCLSp6umMJG8QHgL6u6XknwWNMg2lXWyl64sRp/ZfZfKMlXvr+4t8IST2
PjYehjsXtMG0og0CLlV2E/c5VBu0E1l/mLT6EONB9OAh/LGWnFsMgAwdU15oACVO8jW/1xXUjHba
awLAiBmrZDujHsPFivoV3wq+AUWWvx960VpK2X+q3fi5gb9o95rAmG0blyIlYT81z60/8YHNM6dJ
Nj1j3/wBjb32bhV39Zx//BJnb5PznerQnqBStCvePsnfxwdEyn/jgyAkOaVioV7Gxb/QLnBN4aDK
vdZRQGFc5t/HssVDj3kv3GPbNqxP9gJVdUJXkXNOqTMiwVckqN8cISjvtshwn20hDrXTB6fIvB50
1vXTPgJRt8mrdkJfzWrVSxrBeExfXKSZEInjTbL4JTjuyNqes5N8R1NzS1SDSSYG91+Q79LQWm65
phtrLe9EAoCd1WgsKqxWxKXubLnjL6kDNsRX7VCHWNYS3qHpeCCpFgWnhOrpXaxMn479uAFwpgRU
PM6iZRbWJ9UYSAmyiyn4YFkpl3FAroCu48OfLtVZz7RD/3y5kazlDQwVDrnitroGCW2x8HO7GUha
l7R0Z0rHJbxaD/X1cZDH9RghVAyLurwKluD1hlDIyWyTEOEGEXEcwDKqqG8/8ScPtKSuDgQnmLqI
7ho/jbVMgGKXXvQfwyPX5SNWykkAPr45gXCTHVK6jbY9lhQsX6xFh7dpUZcsNNCQ3wl6qgK4gj/5
WXpUoZw7spt0zYe4ch/wxRzOzYtX5d2sB8Evmv/kBmxA0hMqHAFv13iTqMTPayzNiKtzRwRfEpQA
3TCqDfqI0dbR1av2aIoQZVbp6JZrJu8KZuwWMjxM2tDbY6fgqJ3hskpuI7EfLZmQgzsv9A0zZbw6
dQs9gazXUgtCrqSAKg0A7pnex/FJmho93M7OrpipBXzE3r4U9cbekaIu95E0U7UW0rIO2ztSNgVE
pzr/LIt2PVSt9LxxCiTCBH577samTzywEOAQpMRiM9CnDjLRyPiNHRgyXwf/3SBcfD4KpoWlnPrV
vDVZ000s46Nrhtj3MUFKUPZe0mPuIO7lQFt5P191YsVf8G4x3UbTmFasEwUPI49ApLlv0Im+30jj
8Y2pXqm95tcILyBsbnl92evUKQRaSypO4eLwkOUno7g3VX+Fd2DULYfabvmOBaDtwMKL+pJf81iJ
jKfkHCnu7Xh70CdQURC7s2wLC5WfoPOlLBdGwM31co3BpnpQrjbzDY3ki4frwufsZiKa9s3kYSS0
t3EJdTiMsEPyhK0aR2XWnzyisDj5gLE16BmfOlzSwWmVUhBCDnCMCzM6mqh5yemfKR7Mpz0vr19a
Cmf27Z9yBZig4EQkwsWBWR1quArXDH21qW5VjYTbiTrqULlnw0ypowPJ4kKnjV+QTM3wyhO/FcbM
sUxeH5hMBs9O/vBA3e+vdw3Q8qThHEDOW0o8xMfif5gYpBEbNyfnvJizYXfj6sUrJpeXBoO1x8dz
6LNT0aZIZG4lgsM9EMZYLONS2XzIC4s6PZqq8orWfCU/FcxzZQUCFMam0ja5gMFaeqIIHqQsjeD3
lw7KbxpBSaUjFJsnfLaUoGeOSmigJ1MomluK/U8kx7nsTlki1SuNCp34DXL/beIkv487VQRZBkv9
tVho0E1gHtGiUUTI87KLff/Z/nUjhO+vnYJzDSf7kNx7EwF8Spaol7ZuCjq0Gy1opOVsf7fAyf+9
6AhapSpZptfTPh8a8Z+tZQCE8v3fPkM95nsIYvGLjL0pjszhK9MCzB16XOPtW8gVJ89lysmmjaKW
lov+udOiYqtmk808DZNVBil9wyQ1uGyEQs/J7dcsGwNQ3MSymKjkTQJ3pl92LcdnmESFERyCNHbY
P0IqWOcDHDF7AmtnmiLyWW23My9qG4rhSJ/GGOhG6Ued8QzaTS6xjgJKibyHH91ddyZ8OxsKZEkM
aT3D7EZobWI5uxkbVEMREx3mjx9yVz9QX9oHuo1QEA4ZvqgzTkAyptP+VRg4uUfYoPALZbczLokP
XA5Fto0/aYYxaXVsrLK3/3Oa/oETDt1FWcueaKE2jOLDxslG00GA+usr9qjHszoIRb6oOl4uEltl
4wrx1NhVqJ13bgHO4SiNXLqQrip8yheuwNJJ2YGoQGKErY/tBZWghYUzpP79EA9fgpRKWT5z4be6
U4U5/sPODKhi4Pv9M5F2FIOIlHbic5Nh8olL0BLLDy5bLN0tWzfE3KjcLoESk/4M4tSU6jYNbP8G
pYZYFpC0h5pbZJy6Lb9gpPwXao8XOUMgRPAYj3I8JtxWe36THsJfpxLfRAbY0ogNvWJlGTw9jyml
l7X8zrMo9E4MyzOzrZ7kCY876HQP+66AWe4ObXkbZki+UGO1yU/SwtXughO2TKuVnjmQYGyjiBMM
k/jAHUv5wmFnWNAXS8YGzEeknoRw28oxmhir0OT9ECetp7Ke1A6HIo/ogHKf94eExYL+U4aSK60g
1+/zwBEFlZ1F2wwdOscDQHABQEzZh1sblb84KDcAbNPsPciQVLfYNRbvKRD28U5TMBVyBjySFt4B
xnYVjsgvSxPCW9g6sdjehbYdm3mjBIFo8hwYXj6dTQ47AyEZhgPfd4nuMvqEw71TujSIslvMNBDQ
r642hhm8qXIv02eBr9aiP6DO7uMfAHZeGkNA/wNVKxyWrFX6M8WXJ1Kem/CWASfsPNSsWYD29d1s
74lAASjeRcbsc683HDs0UsBp2R35Rn66R+McK9hcvDv7zIxvuPQy7kbkbx9ltlxowE4pVEVmyGJL
tjlBkhvfu6a1Hm/ySxMNXFNrwX/N/j5Zn8SErrMlxV225swKFs39VUV1DbX4zyeG8mWC2s7O7pTw
RRgr3ISD9CUhYFZehzzHeowc9340rkfh3WqyM/ZgZkxrLWNPc9QR1Eh2kknCoE2lMGNsUWy+VNQu
8jmCjJyKnc1gUMM4lzf59I6UPLojWcIzLdZu/7REXcinkNH2oNeqrxZuyRQfeEhSKJVeBxmzirVW
ELmGbhwD1+UBKPwS96bmR/uTMDrweLhXDa1hKRqVRCPyM5W56b+/1T4p6zMavuGKq/4sg46/I9ik
bS5pesSAtCJYZmZYJXWbiz1oiFlv4K/HJDcrfUSBTgKVPAItVYDO+OvWmHWi86mx8by/lfvxtER+
p3qvd3xnqqcSVAp1s1BCAj3HTV0p4F+PSD229gK8stytNSHxE9upAOIL/XHhrdCRW7Vc1GEpIRAb
H2Mhc7qMPUVwU+s19UHKB2dZXQJghjlMXLWElTuXRYqP0yTIX/JnJYIPWinqhXan3v8xHP5Qcx+d
8cIKUpXqrca9oFl5VH7+TODcnF+mFp8SZ9EPZNyJen/2QWkjZXKOd/I1uYGfyxHrwFWvlAfhYLRo
Fqi0gK9KD5f0IO8myLZFb9AGYUUdNV+BeSUTeZUyKO9O7w7EpgRyhlPhovvP/ZAptGIrMI2xoK9R
89x+bEyBb0rWSov0C0G0mN5rNagI3zR4RyMbwFe0QAw336cZxOEak/vyu188wQZ+3XFwG5lfxJV8
C4C1En5luOAYdn2oW1w2kbO+K4jCEkh2nINQlaenHHRzgV2efgSZf8yYTtZ9irfnXkRq4jSO+CAb
jmAjGvYxGaw4PXPjGTPA3EQADeQoqgSVTwLK5UuA+W9TmmZzBXPiVrZAzZ2PeWoXiHDCtooYNEId
avQtenxp2qEwWH/wHUCFfGkJO7r/h5mJxH6VPTqnF7/PpKgTDs4bwV+FbC7div3h5yF0q0y7C/U4
iaRxc3RINouX8dz4EbbCTUy0fl8kOv54hw3OdZZOkkzBD148rMTID7Z8zcA+0Xz621b5DaDn5Yzy
Md++6YRtHzbW5C8K3XoBYg1/eSlaZ9O8Fl7oymKviJ4k4TxbAvnnwkfwD/bdbrAqg8g08D0TQ09+
LY8MHOgzsoJGPzdQUKr8OttvgNp34Ha2nuBbglKQDSuYJ6wIPcfD/XgPysqozdftc0jzxhfU31sH
BuPHBkPujMArX2Xzro1aKty64aoukuFAKrdnJEPslttGhKDtjz0+ANb/T+JewB1PDszAwmhESYnm
4PZ8vQORSf2rbA4k3zmrFw50LK7GW2bTOe5fSLtC1mBO06LK0U3yDe717XlSOfz6wKCY5kzXbohK
1CBd68WACIr0cAuVkuVTzAwtMILmcPjGbxAh4tuegOstPNchTOs9yIzyoMb2j1oMpaG+f8Nnyly8
l4+wRdrNC1vzVbxx5DIFDq6E0IpPX8g6xP/02WTjhgvAOIp0OIKDdjlVy79xoLeUcM0GIwg0h6C3
LJ20yS0QlP68FibcUrvDQEqREZxgGEOKHB51rXs0FXdSXLiym8PfIoqxuZ6UcZZQBrg1S8Y9lUFn
G4v2lXezfsA4J6VGbj+MVWjaQku0S0tl0JVYBtybrTE3CNOz5GAP8WF0r3BbAFzG58yeVe+nYy/j
zVtgJtDjeV9gfHcf+PtU9KeBq9jFSm6nRn3HttZy2CEKPKJfyt5XhDaVFnRSTiXdyiDqYoif4tMC
lRm4vpyPzeJdaijeFMLn0mYQnxH/tdLwd2Tv19fWCm/kjVT+8KAOR3PnP0wzkHZfyHic55W0Yn2t
sSbcDR2sNkZmDJUvq5a9Sn4adqgOK8EQgKaA9EK4PrypUvkAPPWa9ZfRZ1zfDGQ6UaZYT5xojPw1
nu5MNuwMgREEb6XoOZHtmtaI6tQGuoYzAtEzJLmlS/Cy7Oonb+1K7G2ru0MyITRqFnvg085qe0D2
8aYcL1myfSeYfhcdCXiutpK3Ye6dzCW4lMM2eyrGGR77aCiXLypeU+Nb7e3bWrOG/Y92O7dMH4dX
4NAS/KjjnQdGI6GPAc53xX+FCGtY7fRPpXCqZoWtrsnaSXYKxwmVCdHLL8rWqGKegRV3MphgEoOq
UPTW4IrooYUMHAzArhGBSJeGaWiSb7ABx++Yl/mVXRk+x/E6KIp+uItOr79yZG477HRQvY+KTbCh
4ndJMCo2w/brDdpBI8ubxkE16eDWkIiFRgJ0/uLoRM/Es00vJHO8JKWJH/0Bz9uhDaABY37LI4Bk
mvvgKlLUzwVQqiEVvjBnBzvKKVx8rziRm9e7VGorEl7NT7qipgJ4KBaE4NJpVxZLvCKlp0AiW4uW
XKLnx9Sv8kYzB6FTG4dZ8rxdf0HRsQjx4bmxCf4vzxbsDu9rb8cqBLlEHOvdecOr6OhxgfMJ7VHX
88gRUXAltpu77+s9+WmaQw6HxBeVvBcPTX0UCZeBd99vbwECRRWDdoy4HccUWhLuJZv8eoEyJrlx
dUcOyo0alLH9tt6R8M+stl8Vc80KMk+8A1ORojDfr78aAjo/LGQ8js5QeokNEp7mhgAw/K3aHyOW
8DGWikCTLUU9hzNo58cCIc3C7Opob8Ic2kJIXI9Gg0CZaYUyhK0Q7biXS/7bc5L65BViv+WdnJsb
Ps3dzCTJK0jz7vDdCkg2J8yQQdRX9ccq7jfHBzZP/G4XnBO+gfyrqRiSTo1/5Q6Z9j9BCLDA0umB
pVtQemw7XX6vKy358+nAUlX2tRu3lzGq4K+cY+cVj2h7Y0qLktvgvJ+zEK73qMYHEhZ9VYBYhJQL
q61ci4PVwhrZtm5FGVMZb4/klyOagpvD3edKOnTsFrvbwC2t0gteMXGK7Ip3wEksw2NC1Zrl9VtB
RaUMc3bBy0WBmhcE4q4Cl8ZjtytfR0TMz9Ap7g4wmIx8kNxFlXD3Io+Y9DtlOQTjazf8v1Kswa+0
JVoW91V0Zutq6gXtfddapEugTcPOFtt/jVnHmwP/Fn4l9eSBv7ZZAPL5zb8sH5sHXR9voXsjsA8R
cePsIiby5URkTPd9ph27ZvclxOZ7yw8Hu9gcLSRjgragYBSzoOMprLzCacvxs+cKFYYYCr9Yz3es
EukJsXczk5my78K7iCv6FUvTSgrG8cDwpU5fJEX5ZZ3l5/d1LH/3pzR0uW0x3h5r9acMJEK9gL9X
05LnhgxpPsNCt0xE8Vm7tPOqpT9LOWIp4DFwYqmYuMfSPLWuslrRT7fTgqOdDBYYAsd99ikKJEGj
k+qoSWyVJ8azq6PQnRxUXlZ2cMASvrkArECO29j0LZ+qgrE2/OOeXqq+nD1fDWPoeBiEABAmC9el
Z2xAkOsPWkPrKzb/sCMG24/NbqhSB/zS0t7exX/gkxf/TJsVZhRsoANC1onesEaziJNslNCiO6ax
Uw7YgtHyOEX2DwR86aD604pdUIXhVpjesa1fqisatlYlgdWJmTaEK53F0nfQv9ed//WA6glFeiFi
d0F/H8JEvmF49MgSqPt80n/Y6bJU6TjEbrEr7ewX+9BdGwnv7wxcPGHmOLh7a9xj8oNX4lqK8XFG
hddJ7TTv8PxaCtgw8G5hzDgIL7svx2yuR0GRzl8c0kD56UXThffQpVUO7cqMjYCjwiWaRsPb9zzZ
XQ2gmKSez+nncaQwRPD+jQKs4l+wnzbA2CX+J06docjs/2AfXtAWCQQesinnmGyJINEWiSxAHLQ2
dAKy2DRuNyXlzBtNOAt6EDKVHXtSZfZpqJrhuw9RZSfnvZZpWdCWPW66FGjOCsGGUuiHBvUHvFdm
qRAEJfKZTH3w5YDA/q7Usi6cnFIf2N54aKREnCtYpNCxq9AewuI9WY+YkfBcHrptzZi/XCPVz/HG
rLkBs2RVcJM4G7wbm1OXaANWVZvhTNc+yj5Z+4I8aIi1Yb6D05Uky+F+h3u09pzJM00ItfPkSXKc
DIZoqT0qzEwTcSRx9t3hu7UVwGJET9SOGAF4RDD7oDW7IEQm3pBTDM03dG2ulp6CvjRlrFxGAH+Z
KAZqVUEcDIoXIwNARRx4v7x1RohiLPEL4OAe2ok3T2D11fuKpPS/wpWm0YBqfpZyr5ZzYyK+6bzH
9+ut6BukZbqCrBQvfYeC8eq1qC6MGsmZ2gxN7XHIKAb005mMQisrRIyKL/FqZT7RYBLlShJysyad
rF4fHrHgjHZWCgDsnIcs9g8oLQO+dOw7Y7Z87W4tnvnuur3TR7S3AN5GumYQ2T+Yg14I4rY0xIlb
d0/LmMzV9RJxiWmLTe0s4RelmHcQ848DkuQcQJsHU/YDdiQdZbJAx+FX1thU5Hx+HCBzmOFUza5T
SMcuiG2d1C4Wd05l8p4Ssc5zRfQVe52/INhjEnte6ybsQG01v4zstu9bAEbcxJOVYP2+CLkfMqHX
YfXnq4W8cdva8BbWEtqls3nHRFH8fi7UDJUT6suIkEwSil4JkYWYE3XaTptzw2J+UpfhmDXi83ws
6KtsDaYxLOmdx4P+nEA9CcI7VnipmZRZ8/PIGmg1x2ybzBuq2zcKuCD43xIb+XMNtBhV715XuySv
Eb7W+OiLwpGr5O4/VIwrhcJ3kjRuzSQz/pC9QmwrwMJcS8wsSz1/vkmHSYLMheObRXv3iibhhMku
s1WjDjcb3hczU+c1wh3UFkBYjAFQDNgxKci/3xATjqILwlXFuez7TY9gnFTV+QCfAQgnh9hOS7QZ
rFPDnGUp0TQkFZ28oDRXUyJhxDKAkqdN7JgOxrgu2NkbiiH7yl5dT+oU3xqvW9gDsiKhI8WgSA6G
0gD3g/hP45vK/idQrIlG+yow/0Ejr/iL+IOYiv1iC5uu4joNkpyqF4JDdp6tMLTdjIRT7RAgt/gT
9J9rJQUC8giM9HHM308CZLvXLQ3fN8x158esORrB7WYtfvQ1oNU65+QBrbhZf8Yh7x7uhcmCgrPR
HywD3By8ADgYdKuyVmT7JvWuvb2KaZFXIqT0B0pLSCySWUi88vLtCvYkHLB+s3Fcj3u82lwqQnnS
pURWeKZ7CSWyv8eUnjuF7ez4OD8RsLcYMPuw8Jny1l4jrljlhdQqBH/7wbzgE//m/HWVLxhCPiGp
bSRuXD3aFTemVduVkhvi3FwUqQknG/eDG4ri5cAG0Pq3BDtpaP5D1+bRqoLlaKGzuZHJ6rRlxcE4
fYotRaJCFmPyK1h73mG7tnYMY+2aBW83uS6HMWBB6jny95eLUpEqGnni70gs2MEOZPGsDUlrnqoa
YYlBj2gssqtEPYQxUtsKR3LaynP4Bvb8OpzcizLSGa7cLI3MafWt8gZNPbSounEYprKs4QGvrqHu
ghBPxX1RgJhS4a+Q+O1BMqNxa+yC07OEktYag6/8dmOerHR43LCCMVi7euKbNk+NIS77cx0xIiBk
zMqeQ7utwA+x5SXePwpK8D2wIWPKS1gM+CYvhb1iUIUFwlBfvUBRsaVz+Ve4r2wF7zygJ9yjlHlC
rNGQrqwiR6pdNcfpd253oS53MiU2dUQz8R4xVscNLFwySUv6QnKfzP98XVHJvKmA/LYsh4SosyGG
HHMRfIbvgiygRyOg4V/AqioUNow/GhZpq2gfwM7VoVXMAsdHZySmEKOybKbOlwpJu9xfp+VA27Cm
OMbPBO+EQEfVUrx3sGb97L7LAuUc9TP0D2VhP7+vW4w7jJ0e9oQoj2LrNYgxqvZihqbYw9nHuejF
b/PByDGUud9VQscG/bq3Z6N0z6Spiu+dcH1yIYg0sjiZUCNExx0xDtS+EobGU441Or6XL3az8IPC
4NzzbQxAXaxKQlMWI4dOt6SNp8nJppyJS+To9TNd90RuYKe+ybOL05ccxf9b51nnog2sr+ZGeu1Y
UxD40EAVjBvIHr1laZg0vSDShLekYTdeapo2BghNzPVs4xeFiGVoT7zu/fepECVYtrHUFp18ZOGO
M154HqROfWcUyeQRIL9rvH1eBpAoJB89DV9VAkgRyM8yABNfp+mH17uQ0OmXoyTl67gfJibRK6O4
eMzg9weDLd14ulEVROrf1+qXr0JFQ6qvBETR0+YmdabWIiGfm2sVMu7BKjOgVYM4RLYCh8WnIrHD
jWIsjuVIX3yjtO1n6mlgsHLD2tilM9M+4KKNPc+NyjP5dyanxLGrt5f0kF19pya9vMv4o6ETL+/z
Qqib81jAuyrveaUhZeZQuZyfXF+sV2sjOvtW5nyFCKlfoEXdESC4Sv7H1Chzqj7jVfLAkDvqWy4z
jwbiVJBosE9EFQxgKh2zT4Z2kURh2cORojTe8UMt7U1eYyNb80N8UmSd2PPbgFyyWnG4uWOSDEii
OycrWK8/XBVM1506Y3px8Tp2x9Pods/zF3gHYC/XoannSLwesUIk64gedeP159j1SJ6q1UUj/ZEf
xW03clLmKocE/TZfvg8JvRXRZHyvhZve5JE7CU07M3m0/HmddCmX3ZTdtegQcG5D36ATeW3Th8gT
2a5Zo6kZURxSr/ijoBXKOWDLoepVRdMOs0jEcRrKtTCYpFD+qCRyCQaHAVz6M/8kp9tc59cr2iYh
Y2VZBJ1QeCwmStLXT4Z6GOisshC7pqp8ooGzUYdXwckfvYKYP4KNFu28MhGOtAIxph6tnUo42UiM
jwR2M8et5c/4ran+nw6aXLwefJJokg40MNZYTDgUgU9DsOicRAwItpcg8pThquqNFsTjDgvNtaw1
URcY+BDWvCa1HS2kmnbjqMJSzHRbxUP30FUTeTF+jm4FcafQRWgpvr5Zb45x307aMyFFjeNmAkiK
8mMcWz62oCsw6qDyg6zhbahx4EnJ9SUHapgxDhIy4K9ra3ijXOMs8FlDV6J8kJY9d/MlhmP8u88k
Mttvl4L5dXK862cvk470FE2ANewcA5N3RS3iZbeKGVMgPR50KaQcYPBnuKzIi0bS2zdzyQ2Gmi+R
G1sR+1BSacov8MFJVOCUDPq1yoykSoLAdHxtm9/cawm5daIDZa+OHZ2wypnIquDBSQa+OUip9654
g8ss7eXlmejyxxazbN966pOIOUif/ShlHWOWfYXANattG4BcSHXNPbyUCRVaGkoRUSprD2izfxei
JTik7PWHKHj3n0p5VSzgCvKe5ZUs4J2LXDSqGkcUXGmq7zi0Xie18K/deXh1nqgOEhxtNWY2RJ7b
tKSxXGdn7iK1hQkmlYypQhX6Nn0qNby2ULsN+85zFWvQAzzDvf0f9KQCiMymx4jI8SDkKktvsqK7
spMiiO9sOA+6OECqlQ+2FDJ75z5UYRKutp4ZOfPhq+cKxoQgfBx/57ETrQM+Oe6CWULXTt+zMTRQ
PeXZJYh5YHUu9v8ktCtrQtqU3zB/hicKz1sqoxRthHuI862j8IVM28issrFYN9exbDGuFj31T/Ge
BQyEjT0HCz1gM0dVDerkleJTAgL2Egv23DbuCPNQvgQYdq4tskdPVpAno3a+uzKpHCysTQ+Ffc6l
AnqhhyjpZpPg3W0lrS/vIHCBbCQINMVSvBkCq6buOwRsvAyYAU8SdhFG7SwwMXU23FlQXqK0Lr6/
72fkaaxD3N//oAsElWdQzbbzNpv7iREAb3twhqKpGMeb3eyE54gFT5CNsdcy6KNE61n0vpxcjOhk
5RULHyXPinmKpKbiTFETyFUzER6RccfUdzCYEZVsT7QS6S7YlBLYQF53NBLPiPjBM1d/4L8m6HZ/
KysM4fyeQ2W3fyzJkDdSr+yrHrxQOvZEn2hgJd7k1HuvMJW/EC7FIiHJ9a2L9Kyt9vq8GNCMPJwv
7/K9eB0wv/Y1079+Hsn5jS38huzXEkrdZHbYJeSw4rlgbXOTgendhVQ7YcqKaOIQgSJVHduC/ETK
nSF4P/GHz6PNzib1M1V8VQ8gGP7moZxYJN3IacQztyTdxk000lLaPWgEjTefVnhWSNx+nPAqE5o8
C2dxK6LRGS8817Hozz6+PGBB/R2aJk0qDfdFnBjN1hpFMv7i9yIHehvIy6iB9DakJbchIMgNPGpk
6Jz5xTBQ8xf/n6tvj+8f0pTSH1lhYkjkRnmD23xsvyMDr00in/sMPWAjbazPL2kVwq97tSRGuKiW
UWBY9yXN05w1U1cSrupta8Jx8/2LXtzb2o6iSua+PLK3s6vsMZsdooMDR0sGpRr6pG/wg5SusH9+
r/ab2K/a6JLFIPbuEerHXAA6daTwKSG25mheLm+GUdkKyw9UNBOw4kptiboyhYM5hBwQRTEwg8Mh
4S1IzFY9rc6kxAuKunXny9mjBq9QSKa89NCs0iDCM5nLf6RZQQc5HOmfwsAM5vLIt6Gpqqwz9HMK
I0bFMHzmN/OmanpS8PC8M5SiiGmcIw91SCncJu86KUOCcTQ9akiPn/MoHWXJD6OCzWFMysB15aNa
Jn1XISDhwCdcAQnInZEOwL3hiURRM/P3/x+mayAuRVIKMzrzNvCYgBfl54VbXRGo1Vkh9yVZinyA
UBfDkZVKYBbNgMwr6MgLCNZQqbO9/HgbrtVmVfKwxGTcwY0Qu/N8vAKy9Z/Fdb8TJ4/S0qNOqEo5
M34OqjerygilXxzz4x8oGqEtSxuuwAZ1QPNh20jl9lpVBEduhmIoq8/47d9hnvbzIWKATUfeReJ6
3VdwK5PkDVcVFWabA/cetaC5LV0Iwz9JsEqwqwCXPdw+WbcWGztNarAySE2WY7aHLSeBZL+egmfH
OFmTvaiRqRdAJmQAeQ5KKB/UiCgJg/YYF7x6Cs93pv2v2TpSVxi9t1BGZqdE7B7lFMC/5v77T7+D
sOKkIVe4Q966xe5OvfnxiNrAznDPDl1X7TQzGtn1UHvi/sra5XnEAm7Rhbrx5EMPJfNmYisd3MY7
3DQgGmG8TxSihYz9MJNlJUuZzkcA35U63mOORM0RmTRmPR6h76AH3ZoIfki/O33YU6d4zcN+MCnf
o7a6dS81qUsgHwz8wOs3yor+Z7HvKlZ3RX/swcD8IKE1YhKvcIOYmiUx8jaLMPADDBd397D6+s6J
H+IIoKK5qAPwsc10fZOW9zZSfni4SbnmCNFnzfNcDFz9Lgqz5IQI59WBO4Rcx3bLHbwL9eBZupIa
qEmSnXqICcGiWEa+f9XSxU+Jl5NWHYSChUPuJkTPUHi+gInmj6upFfBod1gazIBQTV7dp4cBgXtG
zW23ujME3y4jsb5ad1XoVe1ey5qW1x1Ll8KQnpmVr1lp1ZBqy1Smk4GO/qQ/aSotOkwj03ztimB1
fYtxRCNiy3mqAO9d2hlmZ6wtJFOOO7BgngeC0ycWpjqWfNLvQgiUel5zL7ZZdCaLXrI/qf8AVtzf
t8UD6LdXe9JJ8ohnApPApOmAhYI+vC/c8OAZ3o8YrmOG8Usaqdankp5BxUL+0/dXiFbcxTPSnnhb
2VmezG7ZHxm1Sn6XuPWUI1j2kWPWPMWghDQne93gJz544ZDDp4KZXehhOGbnAAslVw3i4q/TkpHN
Ob1cg+lQ9d+R3yVkO2i7Y4Pjl4B/vvbJR02xWx2+YBiA6949kyVW903cvUsdRr7FCnUPH1IAo2aU
aXA+SPfKFo2WA1zj9vRTwEn4gNjNus3q/lnTNIrvBhve/emY8fxFCaPx/z7iISqxeGHa+yAqme4d
dravWyzMIQ+nR3SbnQDKlbcjI9Kg9Y6MB+Z7h4c8JBBuvsbqAXXsXpIKxA5FJf5dLKSLlr02m7WZ
9/XbsgUs0M75CF0XchME6B1MjwW5nfXV9bJSalaeXMS/YGl0IqJuuFx4BeXPDUpAVTQdzyo53wPl
NiHS1S0X0LFE/2dzTJu8qanNXjdO/sY5wI0fqix4QUtAqRUOXbp/aGNEV9Lx1aE3UkeHpfUJ1SV1
IV1ZfpvJZ/oZn6jXqZ9syBFRCGGmHhtwov3GnPp3fGiJPk6NP31pakbVQlrXgwzxABpmKfOlfF9m
agrJVfZp0WdTjG+TApNaqwrrFuDIjtIrny2jZZ5pu4h1gBi3ttr9YehHZLddvpvpyXCGnntjmMPW
VA7qQMTzLAV9uau0lWufeiTgI/vXNHWeq7QlVfmov8ST5SsdTPbJAPpDk0+Ekm4+Uz8duBJDxsDt
b11uUDSmNenrBvVRATTzg03l5+CnGflhWwrpSZ3V8DP3kMZG6/UBhsNJKn9vzDPql8gOA+hIlmWD
jr0Pvl8v6Zvf1IlN70Xit3Ankj06dIXUJKUK5kmqQLiLcrCt8EP6cHb8Yc1P+oivEGFAdO5Q/7Jg
It+Kn7Ut5718RFLBIMHACDzdktKHicw6zAbon2xJkuTbQ9sQJH5Z3SNr7trQW5vxbxW7FgpI5H/f
s7XQlXk2IEbWmgI3yyQJPmU4UXlSaSpArlYNS6ddKX4l5xa3TQwwFFo13yBD6RBeiR6q9L0lAQM3
00K9s/79OD2gtbgMrRt3uuYb5+QU7iqkdNfiXntjS+30c4RuFxeJUq8KtJgNpr4nc2e64phEvZip
qWQf/++zd6Dn22fy2etfHyIh13x+cRqP7vVu3xUXI/zZwspWR8z7fTiYS2AnGHaf6sA4wyXfomAw
i6ApH+Kryj3f9Maba/7RmGrq2edTrBQxkRNndz04XGprZ7E8fBPqrBOoCky6ryw5qYjJJmO6RKt2
PRqCl+620HjkKVWt7L6JpS+NSFLvsKn2FyjJUoN/0N6uWntZFb5TMOk6dJxBB0Y5gYlKNVqsvHuq
Tv2dGO12tIrcqekgENNk0fbXGWqLDsAX42KlNgZ4BEapIlGnDK4svaE686Dzsm2yILyHK4Mv5VYt
Id8+W6ibKvd+L7Wf2TwR8CM/U1/TYp2b7jFebdTM/P52dRFtXZOPigZ8B1AuT8pkhwPCxzwQeuU/
+KDMn9mNiewILvC7vQZaj7H6g0V0tOJAzibuoZ/fulbQ+orq/iRXNbSxvjRadhqa9q/YFAX/Qbr6
NE4ZVsyII/nnncyDoP53R8TkHeQkgIZ8uU4i0ZrHsP3Jx3fFkbqq3NIkTB0YI3LhH5BvgDRforbo
ahrmBvD99QL9VR/UAedSW+Dj0OfkgEHirIuySHQXPlGMgIfKcvyv64iEmx6MSd2h06BxyBG2esQv
cqewFn2PtH+pCdmFh4ATBmFchfaxmj0W72G5Ct7HYSbEsmGfTaxOaNSMT7BXdi8izgRfwA81SnkZ
5GB8AcmZIUKabwQSqJl0CToNh1JzOHmoU8tU/uRpFAdL7lXDG6w12oslbf/qivu1Bn9+uUlmfkdv
QDRtD+s/Q253C0tQe9nfFNy7YdtqNA1XfMD808dJoYIEVFljRXEFWLFau4vlV3pDCLubtNqFjFn5
73FPVf4afZTwDQ1tzGipUQ0cj87xFAG/so9gPRuVEtI4WQaVNlu+II128h3pIDYfYKhD9x3DcP2/
4dTSRQWGOmz0BtCWhqU/6gsxhve5WtGa4ndPlVMWJfR0YYN9QcUb2+z7otf7s6Ygb+QBOBrZrqoc
6js0z5ZFs8w4YdguJviLT//RwJLBsxFjdY9jsY7PUq2fYUtq/kDE5JJO9kkW4FnGY8/Uh7SoDPSm
N+zUocQsycioz1DMzVZlokwp15hI88i+LDjaNNJnKLPBZFrFMfxOnZyuIZ2eSRxBHmc2rCAKVrSd
QMb8ThMKxrYtH9JC3KN5shGcqp3zjK0TftQ7xpJjzITfwVp26pThqseulX7vFZPOy+URVXeveWJ9
eAbqXM3CA6Pa2z6kyV353XZqrnEFKKda5q98pd53aAdwHF2F6lrHhuSg0lVnC1VOI8D3jnxRxA8y
pkrAlsX/vQ8kcbI1AHRRlRdsEyBCf7Sr9H5PdR0kkOKBfXzsRBukFbd2MGmm2FYGke/pvEdl2SjY
xVRV54lpbeV7RzZThQ+VMvzQz6pHLP2Qtqugjg9J3fPyyERaBpLe0AZIL3zn+FgjsKeBFWRlZ9aR
bw+4np4s8ZmiglNV/LdBg/GSfAgwqjqlnaFT3vejTT7FsbAqIGcKAgwm8vKqDfnu56ysLBFRJ4Ph
1YKNg6qMyT3s+Ek4+djdqT6IkPwUOtN/wJqIyJ4FNLJqtf7HkKxm44MfdqCJo3MH8XhtlVnnYOEF
KGuzv3oF4zUdcig7fN7lSqfRFnOIEGl1QK7uSgwYrA+ZtB94/+GcNL/gpuMKwa1J2iI3MGFav8b9
W+3k3WvI1g5upUKQKg8V3UUd/UndtYOR6sTbwgAfGN2ZizsxRAc7oubf9lvdGj9D9Kn/svRre1LC
kT9FJOzXa65f4Cgoox168CTyff2ncVN7HnG9+lbTs8rkuZurp5U+raI671mXhxcInKP4Yhd4ocCf
m1skkd7f2AYA9vp0zChCww80Ghay8xGc8PdlP7MqUqjYTHOrvyhFRH2mT2hmKAJ1uCbUmUNQql2p
CzgsyJHUekr98DvxzPvVuUES0UWveatY21h6TbzV2Tt0xO1+dX3PSZ7qhy2uF97Lf8WrWSmwMJ7M
Cvzk4DoGNA8Yi+IALzMno9ozuB4HhdUa9H+aAJSmvNyfu3uUr9h4UOawwOU8var+vPuI9kGqy9dl
y+CcXQRVFN6purtH4R52mz/M2JwMUBxMU0H9grJaFtkZbwP1I96kfcuVEfNxjSMbRwJFHG6hQd98
h7nOLi7B13ckbaVoOqltEGUWGwel0dd/OhOBZyvTQwsSp/rHJcvhXRAx6MS303ro6sSCdJxILBSB
lOufxeissHzGKR3OOJ1i/F6xX6e1d+31DQjfh+NDkoTvzibOK1z05c8v9HkIcx2UPDrqMUaTthtv
WLRNlWwDPYJIdfcE6qacO6dl/VgIlRGThvjVjfNG/buDZCy+vChORSkxvf2RCiih2ra79fvsIXK+
roUs/EcIwuySVGn0JH7heE6DrJaDTaqIZ3U66xvHLTKoXv+StYLybZ4b/ZAZJjYYhAkojLJPBIpC
uSy9XGo5Hm5AkVaF3yaRetoM3aXdNaA8cJk+Pu7OiSQGRxIkvdv3hmftQAM0ozKHzeGNdTgJtBfb
fx9ehL1CAOBCcMTJknR8GrxhKjkTI2KHBrFBDXA2qpnzgiJ7Z1tAHn+3+trJY/94CO91BIOAMdsZ
i8aDjWe+k42ZtKUEqNtlUlWOYb+1I3v5kkH1AAynmRDPln/CuLa5bbB4HYYLx8FLcMCyfcyxS1tV
0tH8PPQXqSw9bCY7ALgvpswCsSak3IKgCBlo5VbX1CeHTsQrz4dBZYIdjweKW0VeA8cQBwsDZlU2
GqFNTZg1qNsLP1r44y3oC54vhkWTU7QwPrhwJux7pTHhoPQT17OP7pvnP5VeVXY04VlFRjLYUE91
OqRPA79l8jsvNvcfMAX7rfBhKf7/yEU54ncbv+/9B+lJcxc9uCEqQJE0wk0hXeg9OcF1DSLgOfO/
yBCbfOpOXSR6U8iQ+28SBl3X9G7h9ixL+nvBAmMGddyGiqOnO2ej82ey48Yyhxtx9eW32lF/Sv5N
i1zvHcao/JfSlgWicO64Kwm8/vLSWy8qpgHOf+RJj1aQquk+zlCbdT3ULbE0RvqU7Kb7OGOL68Vz
k5QFWIcrw3aJ59pOKRtUiHoputm6FXC2m5+CxlKFqaPjFJJGpOCeP5qmq5xnMD2BWMQT7p/6bJeV
WqXBkeKj2js+J8c9l0Pxl5Bk44WD/2uXEA2cSdpSN9EQE30jj5WtUYYfAFHrqwsJgA7nKaCK881C
rSll4Bzh5fa9fNiDqhDH7jpswia5vpZEszqlCwNHsvftF6kqCKZvLuBKYt1m5/5DytAwSrbjA9RQ
9rQv+DSYitKViJXT5CU7RjJre8beVhoY21u1EjuPrx6zKV39LDx6bUrT6m8A+stkcV62yst75S8R
DvqDCEPhdnITf0bVpPCwUUFW85Maw/TaavtPZpnA7rdi0MNt9E3gWOi5m4O6inOpf6E0oe+G0ERF
CToTUpK0/COYf8KVeO6aGc7u/lYWK0DLeupYIrIJhxeQ0Trw4Z4cRw2sZATSs5NifWZ2lP9n+B2c
M902bUpAutfHOj4ch5RmP+WXO1euJDo/M7N4J5Zu8j4p3fEn/kJttGr8SzUVziiN6+RYf1K9ra+k
9kdyseJswjyfEP0vjIaUneoOC8w3zuLQIrgwWivJYfhlEF3nAPxtk6/OrVyq7I0uAselVHuDmkZQ
Tk6VsJKsU/HH69mWIiAxFDFBzir40VLc8ctRN+XZz5Ux/EQDjq8X8yLDPGYpx5pHa2iOPjdvP/D0
Sk1VTr+t3nMmRORtzMNgNmRUVVIdvTJctHjWS4AziwmclPKZm7qOfclIWP0B9Xdl5HEXCImqfTLe
e50cf0fvqcFE6rusPno0j2FBAgRfzx4Yv4vI8oX5Bt2E4XQwSJ1k5gsADfa/i0FYsa/JIDDvjmy4
SuGTZZLUi62oNBfXZzpPrPSLRPDYiFBGfHpYDE8cr6A6VpULJUDh2rB8+avuuWNx0ey79dz+uxDg
H6OMZljbdyT7OZHeU3CATXHxLKbx4pq8rQdpGL2BL3qvXsL9CzAZrH4ISv1dSMvGgNHbVpeo1/dJ
ZbjOdFQoFEvj9o2/QEzXLNBfSQicIcmZ4okHTfWfIn7Rh/9BveE52dnfeLw7WAh8Ma0qOvBEsTPL
m59ZPxqVh+B75UZvDKyMCvE5DhniCHt2MgM/FjnWCwEYNALuHDiExzgF+JxyQ8sUji5InHaFxjWn
SvTDwCNnVSkcFrqcRJjqWxbduYu660kOqr0vyskZN4yICL+0t/aUFMEbrBV9pkuEizVaauxD9L9D
+P0RdIe/Jgs48H++9N9jcoHk3/PPEMJ/xtlaH5Y8tHAkPHSURznuRSMlPM4DRWtlW9fwCSdfeyKn
pbr+V8EeemqEvQz6ETbiZskadLkSVbzHhb6eqae1DpztkPlAeFIeHAXKcHaDSqEMPUfmYO9qo6Bh
EzXV4yoW9LixlrmN0HisQUfKbfcaSnCdu3P+X0VVQcHOwR8z7StgoAqo3jeurtQRVkXmeyj2qdc3
tNpj/4VxTedYfO+qbTXzwtQjQDurLUYaTlnbWrmzeWOjpfJRTBotPPjaAB3FxidxXOdnlTJ4iXx2
5budacL937Oorp51XWm4HUXDTINvACZz80t8XbyZ6qBjMPQKCaYNaVE3TpzpMIR6Gblo1ToHByNR
j8pvbdNFs2jPWS6CHHkZEFOwjC7pwvbEWItxJUrzC+x9P9joih4XxDW29lJ0zJg2FdqhZciloqyJ
5nawHGK3i3fYOFzDPJyBoi9Ddfygr7dJBACnVxT4k5G7jAZ3ATjmn/sWm5+ExbFLuAAPq/gLoykA
pe0xNGc/iVe10CQRnGGK4naTSRClLYMDKyrsPCNBdu/p5zfrHnbSYQScFxsVwYc35UoBvGw/oToW
5/TczPIHl8c8W3F3c8g70uiyIR+X2CgK3yJSuZID1fcCTmuPxo7kZXk7yJYzAYDN5F6tFIeEiNnA
W5M6beT3XJd4l1BevGNFPDnO8YHrTSjRDr4I9T71ei4OEOevEc6eA0bC+Vf/+BXAdsVR+DGOFiCu
mVQahxixnuCSHLm7OoqqAeAffIjwDJBXrzfCsOgt2ZLvuxMxHZ7w2A4YzwpcFoHyF5ukAwekCG6u
kBZU596q9/ZfOnqNHxY6X15yxdpfM1io6VRVg4bgqRtk4FDDAn6VXkBCzwdxPexqUcVfYgAvIKYB
q6VmpY+47TkvqOgOGh+X2y5G07k4uzNDABW02AZz9YtIggxnjIclXmNV4pyNDyfM/E0f+MxSiSAY
dD/WVCKGCyaKGhUSMlTHU0IeTjh/+3A/FGGjQ9iqq/MJUs8wO5lOZ6+NTKLVqPClSotQPZLpNNep
IXREJOfZgoBmqXeYwaMzH8UfkW+dDtLrVIj/9b9H0CibClx1L9QLsuogcq4Z8HvtMBH6vfHyw29f
F+ynQ29T2iAqG6KDoi/MXTTF2HRIXPKnWsgS2to9SZGU9gT3y3M9bBM6aT/ePWTWzC/B9JPvcOhR
zsG/LAnenDKTrbc0TxTMUpdyJ3z2LfF3hGPi5X6QErhAdkFb4QAnU/Q4KOHP1aIIZryqid1pV9nT
gmpVP/I0c0Y0qf+TwUhcDGoDl3AStocryaIV3EStosgNTcTZ2bjehEv5+zOf+TC2SobYwzblZ5Ff
fDK2ICfHcrXmz3bJdARPIj7Ty4E5dO/rqdfs5AIvOWnHIyiBca7stLn3OGeZmaJbE7MhCoFBpkm7
q1puVl3wbh5xbA0sBOZjhdpZIGFW9DhL7dq3cWVz5/Ly4JRSApgr2DGMioJpxHFbzpkt6MiurySV
eH2SvefO++/TWsgeTCMvwARVvpLSyxMv8knbfMT6EctP8M9601P8bbXvRzNuCxhD30o876/0AHCe
xhQzdqInxUWfoYBx1MunFuD+Qu3FXuemVb/5WpK5Dt9bEy6nmkAwGursNqC8N1r4lzTJaKFrdSTx
cLWxlq272+wIMJcCMztUhu7T5ORm+PuvMw2BcHYyNQZ1GDx2MiPCorOUOnRT+CH3ZrdIqYlFUPye
VHrjeQ+ol6nAhZxTRJVMm6PgLcurL58oBfDIzmC70iwJr9b2gSqphaqoPMHHuac0nYJ0LuBlB7ya
1fVRDvAwgUnltq+6hCoEBpS5GNpeDZEkWTqWx4RLxmAzi16E4E8IxWUAnRDebWHTvn8JoiFVUx9z
P0AvqmGcmgjgkN+lkVJXpbh2DrYEPlu8U92psG9Wc5f8IB5kqwTf6itqfzaJ/gOpl6XAJ9qH9GTw
YPTsr6/vZ4fd1JMukkrHjy9FgIeeaSh2w8i7mpajZpN9OrIPCR8OmAMTBdDRzZx4SwgBOqCNLWsc
tHbwnb27OLe4HsvfaCSdudiTG8D2/OzMw5AzLnK9xcTQGNJ51byOVmdbytl4yZNNGc40AicMCl7q
ybt3daqgYoPpEcMYYlA8a8sCHP579ZF1xK1e+jzZ6wUtzgWi5JtnNqkV0aIM5nUMuxi9TOKnUYYv
LLmx9LUx2FysZw2onbPDhI4ZlNJY2O+4qs80nGuzKTaUX8MwN3QZ5Vvy3nhfbIgRqIeaUJ59FrrZ
G1bEiYDmgRFWpYkUdmbDjUvTXb58TYvIJ7S0qeTRD38rrChBcBO4LrlaziV5ySh+lRFoqTtNuu7J
zqMFJCyiwTshWFuHdsVFQ/R+mZsHSLvD790NryvTA5IJLQ2U/WzYbsRlK8WSqHH8rW6CpzLQU2a6
0LGidY62Woy9x6+91wT2liIb48JM3x92z/Yd2McyfQCvCUtDrK4vyjsjoxiAdyA1SUjtRcWT5NVK
a1gV3FVT4/93mrJKOUHtQ7gVGOrOTiW3m1L0O1pAAoaKAYFPtaKlXKPMIDkdaFgLM5zWvIXPbG2d
Cxcn46YWP8lodPOo+H3ilF/wjLwPto8xJJ748rgrNImoWULvhJnxX+wpKUXEGhnuuxnjGUDP49mb
24f1nKQZFuDhglSKgs30s+YnKTCdnjvhosCL9tXVrlOnTJpg2959cdi9wk2iDulXSdHV+9jalIu2
lKtOrh4WXHBbizjrf+5S7sYkvhUqX+vUF0Qqn1Puxo3BSSwg7M+9t4u3U74s+ovEL5wNWfVPQdAL
2qhgo8791S1TfUwy9X+Mh/zN5Un+Ag6URpKo/J1XIiMEImP7NtXH2R+2REomVX3iCTXckAeJN2B6
qYiP715hdOxiqAQwScAg+vSIBZLCGSl45X0VJMGJ64vKUP0qoVoLlokmO5kaNx7dqEqoIBk78Nfo
QvIZW3U8MFWaY0TSKamCZPF8NT98yWIeOPeCzl+9rbq1VHIhmi9asRxXp+5F/y3l+AlhSX/6XX8I
B3UYzBRK6Hc5UFdbVm6Jd0DZiKTuLXS/5rd1pw2w6FSlaO757ozzegdkM7wK34Xws/J0cn/aVo4c
w92rkHr1TnCFlzhzJV7erQYVe1fYUxATLj3ynCPy/m9yuJoixXfnYpP3RchLMdv+Aidq6xe+ZheA
oWxEfTqoUb8xN1P7eua1VdsX30/e8LbAm3jT2PkpxjpxNTeDHZBq4QeiyYbYNHxcvkwHzjdIIrFm
IuL0My2uDvJYU5JP6F0fOF+EDoKr75eVOvzVbNeqsu9X1t4L71hFCwy8AVImoCwZ8bcYyNqqQnVh
jA5bOMFXiG2oIG81R6SDwjmQIzrSIsLh5onh6SvOQGmfNebydjAeF0BTQAl8phIoamfTas1Hea4m
TGbBwrN3BCm/1Zyt1/d7NyutucuX59jF8RlP+uWBbC0SacrDhhSJkfQ1YSiy8a8CFmWlovVuPTwg
6XKpRLbIrKfnpaT1UEes5bG3/e7foJWYta2JoctOnuwPMO3YZRR5xk+mDng0xrL5qXpWCGPApvge
h6rEI1qaHmAYIDqRPjfP63Gq9jyWJnNLUHIvNluTwfwP2G8cxpi4SD+nV4L+zGwdZSryj6zrtiZL
o0daZbay2KPgo22wT4z2DVwIMLZZpImu/h97PV7sKCNq1eYDWB0Hq/6Btbq56MjFa0vILjboeMwF
ZMR8W7FCp/+mc5g+Fo2VVFyBgjkpjgVLiFcV9rpzTgQ0Km17FCmVnBCPKvLo4p6li64QbUYXnewU
6BX/BjZ45J6DUZdWST/Wgttc1U14xe56cYODIvwJGKcdc7YD4HMA3UTAdOnDW346fipHr7ZzD4dy
uFECqNS3R73hx5xBIb6xCAlXxbetObyqgoY7kEdwfV42oADgnFO2WnD1PvAeJQY57JBjZyx0HvK3
AFLzL4YhCWCK2V0ICxLl9/cglBkR9YCN/6Jw5xrtbE3ibrzJyNjx7e3Ftc95K0sTejC5S4CALUgm
8rbrMq/Kt6GBEkLVhNgPrCqbynwG/YLt7hYOTol0kLnzwyrgf9qs+j4EAH2hZF2D7OFQPAfJjK2h
3scqucrZ+/sMRFkwvV99HBiRJk7vGMOYFEh17IgPInRzqVxtTEJLZvSUwqFfAjS4SZCl99yJmgW/
9uHzrO/ncwvlx1OC8A8lIxWCghSZDqQcbf5qy1XARNF71PPBcmn0A5GWDHULP3XsEhWI22rHdktL
eZoDyVm7eijGxhomY6ykGK6m+BincUJZFc0bPav0oTGxBSwH530MgsMCKbFp0ykgvv1hOcRvG8V7
eY3HHM76eUKSz81+z4D52cf4kZWLi4hpPxldUiMsWKyaLXejULDAC4MXgGU1D9EkOYo5KuB1XMlN
iOrkO6IAVk574XOqq20JIPfKw/IAL4glHACdmhsUf58UBkxB1T9stcKRUeEnT/8ytGPuPUFp84Hb
38hRXWu02U0uNl4mf1FrBSd1w062Lk+57tqBd0LAYTMOXSBop8Aq1OiOlBSK75Z0v+SBIrV3tVtH
7VYjwyn9pUrqrs8HHxn5iMJzS+pd8SPWHcTZhxcw2D18v7NIj4rOk7Z63TquKvBqruIA5ne0snZK
ORlaF42FIwJx3RfiC+Yp9rJLU41Y3T6IozGlApPH1HA8QASGjKkE0QhS6XXSPr+xpy55rgR8vSmg
wnpeMG0EZtNBHXZOSta9m19mpQoCXHJTM9YBaklaJRVMnrfeVF5/AAus6O3Cpk9RfvKk1QmXtYz/
843X08bydgvEj1XgyUj2jUiWhbsDGeiOT+YGcyyR/80xa+KCanoQ+GMY99cE+M19/1gAGNIinLmO
aUn90ypjCC7tzsZztjlSKm+avbhxlW3BBmo72+1q8bULMqVv5A9g2rE0OIXuelTJN/HUZylnYztc
AaQjR885NeSQfcewzcjh0+MKiSgdCvGsnoUTBz4mxl6Zz/wu3ax6x9/Z5DwZCynYdcc8kS1KTVcr
2wBKRB265Wkx6b26gJb+RhOYNMOsKXN1tud/lYvca3LR9Q90rsn5kUqIMVO49n22zXcnY+T/BSJp
pXllVA6Zs4LI1e0zhmbE4aJXeiSs63JpYy5x1wv9L0yThSy+SQA/op2ZO+p0ultCGyLhqwQvBune
ADwsHHi3XQeJ3QmmIHY4oKZD528RlPNbvX3trnX6Jtv9zQB7bn5ahoVeCXX114N6AT3noalHBJUy
VsB2VXKefMcXUBwDuv+g3NjWOkEYu/qYWeRRzKI1S5f0OjcmztfZ1lUvupUbw40OlLMb6lzdAXAA
keM99Im2cclApaNeAdAaXK0Qw+4m8LbqaIGQypzHYsm/0ZDCLbQXQBGobD9zy//1BGBLmP4u3IQC
MmRacL5b4GSOIAq3myehA95jCc6ftrCRnM5xekqPPSXTlatMaWVGYxH0tg3ObikjrUqtPtGYYrWw
aeUpXu+HQj/z85pulGkwutXnY+DIslcom1u7myEDh1jeLMLDLWwbAVOAxa+KcV1yaaw8Fqj7LsG9
8p//vpi6C2mbhYYihxjhVixfvLwb3hwgAtXs8/lcQC6kTEz/KbrLpsa4w19FfK/bhCHq/XZgp5vA
fpBqtJIT/ezYIlKNlAC7Okpi9HfLDsvLv5WM0JXm0RISwupqAj8SUD8ndkZuBXhm7Z0gTh3yT37B
iNylEtRR2+mjvLHx6WhSqq35BM/fXzwQ791z8Dd0XXRb4kDnOvbeLKN83M7TSsdoQg3uE2XCOpn5
GWofm3Ref6eg24vxP5vAIyxhQFWhGLbTVuf7uTZWJYP1RqTKaDr+9ujkgwjeTZm+p8bEilYhu4KI
sPJPxmYBZI8DfUyrGVOWXXgTz1r3KdclynmCRmHWg8Lw5RSMQEPG3UjmGNN7xMMRaxk/zRWVekW5
R1hSFzAk6HDna8jzkCVnKk0PzLYjn+cZdgdhY76O11a0yIKMgEIYyBQ+GDo6AUcWhvAldvVgvtRK
sf//xIV1TyYZhH77+mi8E8CRB431jC1Ui52ZQfmXpFXlhyWuXdrEXnzoDneMjHU9a3xILRvuJ7vZ
56Dpf3utIh/e+SbGx6taLtq8CM4eRWBFnIHXaQZQBQBA9f5utTf4VZuzevhmJ9XphYjnF+dpm64U
lvAehfmu65hkg5hW70eA/CKzphnVr+gR2Plp0bmcofba7RFOrBrJhgLxK3T52eH7HrkJ8mg4l0SJ
TnMs/43a07pq/p7QsGrt72q61+qkTLW5IUOt31xmzHY/+JenKyAZsfzlNVxnI/pzomhYbML+KGX1
ymLXyiQ7tmk7uLt67715n+xmqR8JbkHrJQZtqymDrQJQ9WKKOiTVkXVgrWePodZag5UwWRpNTpYa
XwdiCh2aEITIjMutX+qd7Hb1TOx9eMe09NK+Wki5ybbZGiFHtYALn9WAxTEAKOBIkHt3ofsGCOvw
gLnkMkifiiJU6HryW7e94TJVoT8+hsBF5lLK5VRCCYNn1EKcDx1U4QEBEJJmneE0Njm/70mXAG5m
KIM4I0IYa+Kw50nyfUWXUD14YM/S8jOIRxN0DfWfTXqj2Fa94z3I2l1fAZFKdaA8hHGfawPuZMvD
MJ88Gi0vDf/PejpDibwFViIz5TaQQEMbvlCsjce1A0PpYzx1bE4yEVhFTw60k1uc3yGz3UlQfYSf
uP8cjofTKMkn9IS5Veg+7YcBIbCMCOgYrvSX4GE08bOs9qC5+F28oYSwUPXoIPAu7ie0ZNKITCGs
ggoSo/+90odke/zq2e+NhtqPAkFrOhtY6eDVw4JzfFzcLhYAgH0aTtfo8kdao0UG7bsa3lL1rwCI
EGEb4YfsndWvAAlMt2fLJ/QjyT6MqV+Tdhs3AxiOyp9OqhgTvTdUbcar0SoqwK7U3a7TmXSoIhUp
PhlOl9soqHBiOFWT+/MfekKH0rwZDwj90movjNQ+TSKB5abhnsENhLI9jH86QUwHUxbYEDs3vhPn
M+jHs0M3aJyiO3zw1gPG0pkZ0kIYumEekAmQ5S21FdwKq1aDuDfGB/gscRLYn3duLm/75xJLSNLq
tfS00NQ5oxqYLDYQettAku10E90GHrym6+Moqd60+I9/eHkzq3BYn5+oaLHCa7gl/j8K8htvqak0
Xdha18g8nWFLjE2W8gbBNaT4LzTF5p7SpY4hjZh3sglxjjEA1o8KSkpFiyjZzrXBKFyK2vubjafX
82/2Kqdt/nDI0FRD9kWi9flljpOka4tzvZsPbFU/MYCbq/HGffzdxGqTZW5YkJydUX5j9LzLlNRq
ewUgdjlYn5IuAGLh003YkLXqSaJr5S+iUVssAypMfwQiPLQV+2nfW4WdRANFM5vlX0FBnI9PNjx4
4E0hEUNAxeykFYGXKQvS/3yNmHZlnlZMTId0PemMDmmEI25DMkgkWHQLI8bDEDL7rhrpz65/9UI+
q9hVm0eD6EULVa/VgNPh5JDuH4fsjw4J8i2+K5o6l4vR+eB0hSjdJTNKsO9x7YK2+C2IW+F9eyqV
904q0AGMX2/CQOTvp1bOYJ0NIKM55KMpDOhCoIi7T0yhBJ8aiYhI7rrP4SoiEeDwYULwKoYyrOyr
+k2atkEGFg5kBsZM0LqjeCd8o85yFFl4bAajZHyz6fJlVJ//jp/s4lpibpG67Fx2O+o0PuzXPOYQ
T9iN5FivzLYfV24EW6suVY2Oi/6043d56qtpYiinP08ImSRXQbtelt7Zxqz7zDmYFeV7elWSSWpd
p186ri+tgh1SdTXpAynd8ryyEH7d3xe9TrvS6LQHaQ6aiNGLA8cSWRTRu+duVMuuhMFfU3R2b+/V
nBU/NZKpNxlRF4kcWGAXObjGGcw+OQFDSdF8bQiZnZPlwjbHl2esnfBu9De9H8NOzgLnBXNR41RY
FU9TbKAt2qGUEJxmUJpyQ8l7hyU6G5CyNrjhS+NwFJJM7moxEQhQVWz9T7AhHhZorGsX/umAZiMY
UIp3VYRpyGigkHLzVB8UcNaDRH9cPr4O6dm7BJfMX+3vLvje8MZ49bFR0FzQwHNvq1o/2RHSXPce
wd4d+n9hl9ik/bDZnaaYkaFd/FKxk6RGvOQ3MaVFpVtnvckbbgxwxOBV3cuT3Zg+1FCEi4EeRs0T
13ooH/yll4xL3q2QdjFWnn7N8lbzwaYvtEVW5JjWusFfyF7pBZGKvd0AYNWFFHS03gGrpgR5oXPw
LmwNiVzqrPuJ3GPkt4PujkF22SqGwN5FBo2Ga90VG0nrWUB94qUyfiLUgoVpUIkqBrxbQfxbSRWZ
XFHCI4Ct9KheQ9WhmUhydUlSEv/Yk9EmgGiiH6O3DGJCtNGVGJI//0Mfs7r6k8DxVfQMsqFrCgVy
mEM1bK5EFWxJWJJU3Fgd/9jZ8+kOFJ0YvEyZjVHfgXUWNFMA1NKrupY1mLzqP/lXfkWBlATZmiL4
Ejwp6QskMq2WynRyqWifUPgjvjPRkLFmBtFc44DhILLTnvIpyVoB8nFdkCiiJqSdUM8u6CJHfMk3
IZIZ+LksTbYY5xjTg6VoHTWxJrmNadWZLxKn4kvZlwepIJS1ETFO8Ae6edXF89Oo0y8h6SOD7ohf
bMtlJkcRLmqEaUFsu46LYpifyDRfiZszGbcdxgDDaGkI+mrkwCc3elf4mg6vX3DX+rJB6rA1eK0e
P26Fam59ZY3xWHEDoPxV4cgjy8oWEsSfb/ySHMMlRaVVhhs1ruZUWbjSEptKxDmoJhTENhXCfOi4
qRh8xwW56VPvhGnEbfQ0uFnxFAARFftOzVcD4gr5KKwgq8OqdOW/9lCF1lnicljwKcJMUgfckwge
W23/ZK4vZnFURPG79UGS1T2WzlC0+5FAwzcn/FP8YOvPcmwzaTXcLjD2IlWIfj4ciUZTLiAYzAeC
9DlbMKWCHZLSsk3v3+NeyPxT37GgUEI/FC0wtKxHUww9pJ/yWX0gxWNz63Hz5kW6/gf1CT3Rft4N
TftF2vEX3WHlrEAnVUL0+EzHqiVnSfBcRvnkp/mVqAUUsjmej0VjfSEL/B+4jgUNVz8dNy3EXQUr
Y3IWHgICmWOCDFjIw7K19+6SaBqIjLRqDZA3P99xsDSIDoLBFAPpRb6BSKffviUOrbfQI8+qunR8
qVCFAgICNAPpfRan4k1Kzaw/aoAcGCouRbyVCWxCmjGs5gaNsb8oVnMnuKDzP28n2thqrv2xezQc
We4Zs+ix4p3Ah/IBg5Hb62esQ/B/qw2bLJI+zHqmENln9M+SpQZ1orZPPWuBnyQBsAsj98TrUNw/
NOBeVf/P/XNOtA9QwevobIEUmLF5yyV+50vdr3KXdl77nE+S3nfu7iAcv4VLCQ5R+QmLejF8W5PD
YO1QP4zT78avQeTi325/QNGcTRuXptd+NSsVpYfgg3I3ZriSWM1fOV6NWl4ig66Ie4Lsad0RCul9
I/E4KdM1c6o9Rj1krYGbShiOcYQhoL5Enqe/AYDuv6DPtVhxwoCAEAe61crPTdnbq3bGakiZsr56
UQ7Ykc/C0UhEpq2ZohSgI5RnOB9ScaSLznHj5Sc6Yqpb69lozXXlCJaKbrCEtJwWjZwWw/Hhd1pQ
msY7M2xLglJy8rgy1Id9kdofydx1oqgeT4gPRhq61as1Pr+MX7vDeOg0wddWHnWPaOCHtSVAKW0s
TMe6QFlg5id3GM34XzFiMG+gGlKi0JQMfhNy3wjrLz+p3NToyPKyzvLym9UPiUPR/MVKnrK/UWoJ
vRmtC3fnbvPFIv+l9b1hnDnQ0kL4orQlUbobogDb/ZqnJWn246P6RRuoQoLNW/7g4Or2Yp8DNvwn
z4wmQH2tsbDnob8uf0eOp/hG9X+Grxf3+5ZlJdjNk0Km7SXzAlrMes1Y1SRS5lO9Bf2elgD6dpIo
lklIoSh9fpsntbxQzTqMeK6H/7olMJbwEFhSUAX9KCKaelHH2Gv4JFkAKobb8yNEZyx5h4cvcdrJ
2kzfxjmaPLWrEe1vnxQ3+Y0if6Udpg/qXKemvK/rlXSjP6x2y5LJUcxsLiOgujAFNl2KvpDBHKnT
Dh3rxnnRyKBehfm49TajoYatEfG+gKAaImCmIpQDaD6xIfGzTaz9H5U6cE7i+IEtliD8HrxlKn6+
WwCqYQkDb+xOHpEOZ5ockqsyYAQVPS27QoInpB1qk1ry+yqj8ok8S1O2a0YuW5kRLROaWrHuImZv
3eBdh1bv3T8I+b7uiIFzrke3hyz57jAsm4AuuvNwfBD+IKNk6Hb2Vwin4nnL6ikG44yHQP6A0bSW
W/d55iJrIuIE1m3RAjAZNwld4Ig8aU11fpDcXCTHII6mHHKOWt/neOAmxF+Pft/seMAvEzFNnbRV
R5c8ukCuzd7KQSaP3jLcB75p83uHunONMmdlJXL+HBkibBQbzUIkpLFYrff1xVlyOBcnf3tI7Rn6
Mh/LU2dzcxXBuwzBTrqD7XEIGp3qmKLClzwOpXakZHSy5gTlvSnbw47GaM10Cl6Il11Z5F1bKASw
nbWsOyrrBJ8S8XhsaFkW13f0OdDKk/f1nP1Ft+naCyZe56TZ5npQLPRU0FlpxBKtHyoh9iYVi0Rb
Jz9k5v4zDkQmkJquFhVEv0ozCJdJPcZVhBD/DN9vEmFABMUg6QxSL2siHVtiTtTzl7XJ8hmTYHWl
znMKGtd6pbr+5fZijPSFKHC/TRmA0E8qNt8cRP2FhOb8xyrrd17OB987SHIlmgbrpG65UF5XKoMw
qV7U7WT+01/UhMm1Ua0SKn8LovxJtl/o9Gaq/Yd5OxW1qANj0O6lJfSqW5osCadl28nA2DD4/FpY
ynFNHkzwmXoLpqBOtoRGGvhUHTeqVNNEzSfuYD9jsILemYtFPBz8S6sAzHe2crI0XzKh1++Ip+OV
H9SX9Q+r/dm9aYI0aN+wlKPioPSE2autRctg9y0Tj0hz+skRyyd3UpqevhtctJJ7/Dy/J1KVnZG9
iuxe5u6YxZUPMc8cSGg3heCKfDSvhGKxWY7+bMZqPuE0o8PzHb+b+sQPwK20lmQeK1Tg/Zm87B2Q
+vW9LbaFUke1JjRZNhPibCu+OY3wIvXx+j3M/Bc6R9TGF7qcCa0v7lYkR8nUznq8SFRVP4fGIcUH
2xJfijoGy+NhEG0lHs+jGKi+bD2nr2U7VinyTSfpXpiE1dVhpRC0XDAVv/qX0cOF230sz4KxIJOu
/g+vMU5zgE0AoFPD14eL9oNX5UbkBZOWUw9giYK0+SZeT6gFU9VJb//40Al4iohEOUqBAb7EYUng
IwhVNHCTORsWO8c/fH5uF4q6Do7YrgMaEVPKmVqkLs9+96I9/VvYjWTUF18yf9gB821GouLL8HrJ
Jf3rpSofd3jxlx3MnKaglBXSLq4fvoVje38UfpPLYoBAD2DFac5Ao+PJQl6+z6NaUfQFVZYk4wFf
yS2Qg+nk30C4iYgL8zQrWvCizo+pHLq1P3Eo/qZ+asysYAB3efTa6/4jnMZhvIq+aCr1YFbYI0Fu
8K4F3n1eZYJlEuVTwZnnGPCRgr+R/bI/B3Q/UAxA/lMHUlZHHaQeQyU5I3dRhGC2iECrozhHrsOw
R+CLkLdFOoC2k3lAdOtrw82gEOcOEtMTj71DaIxNxi4exZWLaiOzgM+qYCVNHX63PhKTycIvyt2x
Lm1dq4ZwdinWF0AfOpNywwb+0PuYyIqYuAGEPF8wlM97Oax+jNhui7Rcixd2vVTdqOfKG5xYFD+l
ZDGOHJSGHFlZRJzfeYAIHtmjxvG/IMPOVixC8TuIBVxNaAmpvfA9t97dYsp4ploWoAcQXNn0KCpG
OT50dPlEKl+m54EyWnkJTrgrE+q0GeHHaiyxwuCQM8cLvmkeNWO+dXuVnFZTO65wo33F4dXQgr63
AQ0Quxqyk4MKaybAuvqbrhzXDNj8hhitkdhXHkKxq9m+CkWmYEIXzLgC68N90keJzI4/+LCYoNUF
PofQsmEwgIQEBFa+hSJvmmTXOPdgw3Gq2uVBwnxO3TwbRyO4nzzniohnLmSGu1uFdU2bdTIXDG6s
X59ISm0fKWqN4x7dF2ubgIAPmxT8sH3UHumtkCYksjJUNpcRDewVOpG151YnTixPfXH4YaZtuCah
n87NiDQmZKRY0fRWn1aE9qrcNLuN1q8ivGGqy0wOpv/2HwqiETT7wbUEeQ3A+mOB+ercrVNyZguT
KUFMMKbh6uTkPfutC/HEXGQ3RKDAsClsiAE3D9XfVKGgcugOqeezXIZ7YVf9XWSKYYHSXd1f8oF4
qPsqyEpxxycZkOj7DUIhIPIQ5Led+LLZETr7FhSF6+dFR6N/VF237Q445L754biwVRyty6DNJZ/F
LhJeuVzYU0iumLr3mMU9AaDyOJL1yfDs/j7C/yu7NZVqH/KeMWKQU9p5GgsVUz/Sbdc73E3x8MVi
MoOQsPEk3wlMiDlrdnnzgZ03zPBnn5mGnEGj0gPVAdmaBzvGtKjLim00GynQlaIJnqwASxCyBHUc
wV2xUn7Op7cqhFyy9nAuyVnEuhR2rpt50bzdHQZqViwr5xVdwf7Tusf08xiW+ynlklENq1dFM0xB
tXWbmgPYjCkFHqrALhKm4/eIb3TZrFeWrVFRWpEqs9ts4E6EvjSLcTWccqzknwXzrWmzrCfG7juX
nkjTPrSCCHZVc0uOCpQUiR20Pgp06w8zof4JGk4UiKj6Tz4SMaL9kbr+b67Y+ltm8ZXxQmccu9jC
u6O4FBtM3kGQp812CJ70nXh6E6pncjFuna5tPiMSaUM0EaACBzGdpm73xDiy5K9f7BH54WoauQEu
Gx3G5W65mMUNJnuFMqzNDMnHHM85hv8mL6Pkxtm4sIPfH76Xa1QxlFygxT6UE4Lq1KKonurIz41R
U5FJJvErHv11gPX3ZjAoEB9UbvRGgJRuIu8zJUtrlTU+YAZ62EsMRi3TtXBrtO/NzhsFsUG8RSZB
scJYnZ24d+0CffGOQ3qgPIjKpygOuy+avAll5TOggjoWZvDrL9Dl6+IwXbeQTl59Jy1shtgQwZUm
B7kHoO5DJsIeVEZMDhURNJ6UOD7cqwPSP9r9YLgD3VsDvPqOIibTzAp28aotSpwVXipF9VbfaQZK
vWxAuwvffD3KuZlQ5eRb9DWzVbfuhyoCd+nbh5ZZIKD/sEGHIRRIhmyGk0Zb4A8sp0DEerOJaj5d
huEVsSz4Inqu3cCZzHdSGLz+GlcPXsVp30V5veQPsLkTFN/S+QAbGgayk2kBjrtPZsv0dr186wef
OBaSrG6eAERUNhBTEM1S+Ywph3en633ikP+sPxZfoY/Nm5NdzW2b/D0FIohGmahMPrN3PXZc2YI0
Bk7OyIJptHB+YmOSM8dSUqKaG8Pd3pFLUs9GPOMn7AoP0TYpwOruepRjPrAYJ/gIZBv+iuVoTMGw
6LlUvfuz+gjrrz5qbIUqMZOKMki4frEJ4daxN0cxgUBbH+pJJXZOuQ0K6iGp9PbpDNlVM9+aSh03
GZnXU7PWenqKIJv9ZiPxT4BQH9OjY/BWZQIsCq+Bs8u9DjKy9zwWT5yQYOXFky8Kv9oMSd5+jsTp
uQshccBQLEEeubu5cQvgp+GXbRlDJ32S7pPGsg8MbWf2sje+Cprz1nz6HbcncLj43Xtn1ukREXD/
M0fzfQ74KkbN9nVRVXZzH2HdlViCq75vdP/4LEbG0vSx037OSEhjP15ZDl4BZ21drJDS8NwSvLwL
uy7+JwHySQI5E+Xs44iaUdPVn4j2i7nLI0mnbYInTCeZEHtlEqHPlahVmE/LLfM53Wq/KREPH9T/
WD/HmeNMIz9/1Ksp0sspOX5N3bDDe3xyRSebL/QldbP9QqzR71K3IKCdKotSgdBns50WRXGaUmn6
GA8I3nKVyoDhYIb7XsGyuw+35NOt894251LNzr5t89pZrqCJ8Cko59YziPjYdF/4piB1wOFptOqo
0/JDjPYRVb2vR+mVFFWSu9V4eyiX5Err52JMe2avdUI+UokOarvx7D2xh2BcWNfMMDu2uZPDNXeY
Ku5hgBsCRt8E9wM5rJtcegKLiwUWdq/K9tjXcPxFd3/utfnieiTnXoLYrszlzIMUs2os3ug9SbIt
I3Dk6QuLJHfjSROtiP2PX1bTCh0+Vk+8ARYQozKuP+fRmUZw6bMqrAGbFvjDvLQNNW9MsqrcCq8f
Bjc2awldq/ndXXSv29+E+yKr8Vxpo6vfMESxhNKD+UIHX1c+p0SOEZbXyql3Um26AWK9Z++jIWsJ
DElNXV7hJm8khDRnkmdUwtdEPYwLoVISK+SF5p16iK0VWiwB2Wh9Bu4I42dD8YWkrxdBVpQoAnbY
/L1VrrNFwMDxjb8+oDbUGdIZkVW6WCYk4QeJ5eGVuSAtYuccfO4NGDgdRVtQmQ1yaNh5VWoZlo9G
yFUpPooJOO+7t0Vjb8vPqvwsFq/N9tDhg3TS5KCZ0AtuGQY91oyXdk/F948qZ7woownJx3/e/1Im
l6whR72bXZJk47xkVJ8R6KUaHLXZWQy7o5GD5iFkrrEXISoChxwbjs1GgjrEDIDKkjnyS9it+sX7
wLkdZh1tnVfRC0BPAAKEn/mM54a6BMZSKBWw4mM3tMl+7iIU1ZaKCFymCyLJHPysc4DCdphtpcPP
sEhIdhUVJo0KOB90OmKGmfl97GKBzVfynMjyAWdJRogamAm1YDIm5fH/FTBr/PdgpSQSGjT3Qpug
iipnE9BEotjqq3q5MG7qdwtXU7lLwAiP1O08PqhHip51zcpewP/WW6SA4Hcp23yalWyHZ6b4MXj7
U/nzrt85HS0G/BvGM7R2inJJZ40ThkAsDeIUbWWQVB1PrI/b5xjzTOjngDHw92/Ix9NIQDt7vAlR
luouOITs1nAxDDQpzXlm4suFHU6QMCjXBJUEvFCLMxeqm2R/I/jwmVnkfKEqyIYpuk7hk5usiB83
zlPLSdLm9bIZOuJsVBLNrajXnwfDMX4YBycESs4PLA51uB/+gHuCEHbEcZy4rl7N/RQNmYJk3paN
65QOFA3hy798LGDRM/FEeE8YXmmZcymzAoZvzNiixXRY8mxfpwv3FIzpaEGhmqsLRnWrbQRxlkgw
LRR3tzdy9anl5eWUA8ZwBoB7oLH38YR++arRnchjJqUEQ9ADnGiNWuNodsZ2DneibWivrFXepLu7
8P/c5biczQVdXnNw6gydg/1Rdlaz5RBpbqmLS99O6F0CkfjCXX3o3N6pUnO1IPBCBGKjUppLWbrN
X/6yqH8pVa1YEOw55ovtVEt/0/2JL/whUFpDtC0Fi856w82ba5doStA/IKajmUcnBoNUzTyPPzIV
SOSd30vsAEe6thhEx7HgriWSL+aL0033cAJt1mTskS87GK7ABhporpzYUZ+AA0UWm9uwuiJYluVj
h37eJmOWcI+keULeuqVjGv8Fp14EpKb+2OjQqaW7IrkMl1txe64U4ay14p1R60RHdexcYJEBrl1t
z/1zgVqBVHc0v9OJeBhboKwK7u5BuPsq2IUxyUsGPwNPLq27kIuzQm4Vo/66LMgmhNQfjfeeboN3
WMZhx7SSl3J9raUMlRtCTa5yousebhxyYupYOljHQ+3+VtSTIH3iEhGc0R3Rv7veM1GtS58WlH4P
jlAN994mH8DnTsAWgv0LCNUigRy/q3E14LC9gOZx52mSRDHXPcFnGSgkDGee5RytKNzDQ92NEwUe
Lf6weGAsWcIluX//AfkSMwjFE2PRM3uDp+34GEB3glxDCKXDIyOmGuQeeerXjYrl+QfTbhBCf98j
4JqVrElmc4/HQBX9S5OxVCZigcCszQa2vY9BTkA6z/twK0aTvsnxVmvkHZwo/S2P2bSHClbN7Z8k
c50M6gtTl8RcdAwIOuEhxEkbeIT77Sv2nYJT9ZpvFd04CVi7ot5LFoz8GpwR/YF9DkDAMGKunxkc
W6XukUa9DQEGBRh9iIFHtC+VpaP4gG/rPO0smXKD1sa2Bu88VRYDwu8nhEtjHXF99nmYqXdSado4
HBje7tk1AktHYXvHu1Bn/Qd0dA+1wrtIIdmSHtKEO5HAvaP0j4UprompN2pR9fhWX03nR6KEAfMP
9v0yFP7HGJwDvNZ7etLElnAHy8AAi4UKWjfesmN8pSdxLFN/rw1Uhwp6g4AuHAZNXYDQeJFmdii0
EMAEBM3X5Iv76uo7UDg3SlTSpkob7qRsiKenUew8AXHC+hEPbQ+VGQZtCwKrrHV/oZLK/8xu6ulO
21g+tyFBG88VkMdyu1S6Q0AYa5plxhnHSsiy+O7isA9VVgtF8OSMaxTwaOCSEaaESfa7HLYwoc8W
+RDEXCpllqLG9i26VOIYk7CG4CFeQkEMVqzX7qrWcHuOWBy2BqgAAdVL2BhEU+GvUtmzS8EoAd45
lAJiGtVhd0fWaf7SaU51qAxr+4Q9N2iRlUZd7UXMr14m4NpPNKw86YRYm8wI+s9CvOQE/CbZOHww
pmUu+9BUPU7TQNhGyjzKdGBFTqkkCSjzQil2zBPlxrgGDtp38yFjb1dOMcc5OQLiRBhD2dkkpuEr
PWjmOyuqxXxzD4N2Ac2ccJcyp8TvbIzYor2IZoyG6L8GDSXDLyp9NjG0o9RDr1Wl2bmo8vexqy/E
GekPJvhIlVbhMFSehEzYk1eSepzkZ0oCakr44BH2E9uYp9QF8ewJcItL2vqT2XAvsuWCqv0hgkOK
pY31nmlhzYl1Y6gWgtMFOpcejWNuNjDiufHWkgJWgKcP83ABK7kpf7RclSeIgzsflaeasgmjMa7a
EUgNhcWJCTgyLaUN/MvlgoNmaoiH8Yr0/FlBegwm3rudN0x7MgVTAuUSkrWqUPWp/A8LTirFl33h
lgEzVzjX8Jt04IJ2nQc6ZeMAJKwQ3Gs2NRSzzpq2biodCZe3/azmTmyEo8dPRUcb69S2u/6E+vAP
LsdFIjNF0f1k1O64Y/ML/aAe67ILXon/PeBsfkFFbd7K2tM84lkVfD5C1RO+DCUOa2sDgOoFsP5K
xhJfODLfDTCXhisIm8E8AdZl8xN0N6TmKRHrk1ZNueHnId97d62GiJ+ekLRJOgBcJRqd3moFcw5+
R2djiYtNED40S2UyZYM6jSKJPOP+Qz8HFhVYy8h7bb/XxYDLr8TG47Upo83kA63qBErs3+EBAMIu
f0c3oG2MEyVXiQOto9yTnKBU40XnOkSbKRiEXiLVd6qTWGPRz22rHUMOaTdnKzfcKG+4vd1eWBxE
Xks6apvtHYTdLUDqIs5wQ0CpcH+71wCSZ4QnSyXx98wklGJDVnvZg7xMIq+QNVe5+ETUdonxH1rb
KAA8Nnx+TqRhDK1KeEOV/YghcFR07PVstm/XwA020Hp0BevWhc66tdSpi8UiVcjjz+Zf0Zma7cbL
e74QpDK4/vn5bs1wvHwbLVLcWa/QC9ykmtM3aMJ9qySJPts+Z9dw4pAdpnxhp7qXtjucgPp9KXu8
kFGs2gfMqV98bkSbgvR6KRMNBpvgHVKU+DVHe+IT8EaZGNzaWXrlV7q7bbnTjZolYWDGWO4gzhXS
nGCDG9yL/TQFelJ28D/ZGYQAS7Jph3vDpy/aiP5jJdJB2K2Os9jbnMEjPa1MDrJAykACGPhE54Ci
54gADvmRdvj4rSKCaKOPOTlxFCsfeFQ5h+m4eogAGgsTHc5L23+vDeIPEjiJeUuZyPG2JokN51qn
doYNy2rCCLLPWDNv/M29isSb1/WkENcWnli/vmqxPQsVNDYZ3m2LMwklEp/gcBMd2zUPZqkwzCEP
gPXdhNUQS4Iw0Wr1GIBFOL8IFGdObpOCysES7juhxlpamRNumv5GWWDV4gZQ5mdL4GCLz709ZUjK
YvsBe2Os3Z9M8NHfPzWOBje3YgHND/7L990JvYPepblrO9etPKJn7x6qEEWb/tCQHILyh8JnDUUM
4tIirMJpP1sPPy4v8MlRSV4MVK6jp6ymi2SK+f8Rvlu1oJJ9Y/vc3imAxGQEV0VTmPGR7OdfHW+i
CX7zigTZWqX4UfMGdRsISSau1OPpy9R1txUsrVdsilT/J+9wR8av+WMy5m6OETqCSfDknhWY3gbV
QzS9eIPvvC5zpTmaCKjBDDODLAqy5I8WMmfOsMQgzH2+2uKt3KCmaZb+YhPYzkmITzOTJC/1Xb52
Ep7qF+4RzA989NnesiICrJesF6Qslv3ZwE7nKTUzr/dZMaglhxt4NUyOvetA/zLB3UmrHctQBvob
pJhlJTyfuD09nS1X5kQi45hUY7y6l5ZVt0srQwSog/TRRxINiqxkqyvnwQCZXLxmD09gjkIeElAj
ifcoFvK4zMa7QBZ5XAOHU1vIJ2MyjwKg9F0L4Yi9mEfQu9kvcPV02B2JRgPiWHh+dC/v/a2O4cZS
yuEXx0A/CNoHi5hpZqaOscXI769mIp2XrtC0+wJ39RvkCPcV2p3YNIi/RPlGcsQ+xTO7vAHKpvxe
tGmMUO2kzuEYfygR3qS4Z/661fYrrlHt2Wwpk028+gcYWsSJNyJFKf08/4gSrmujuK1IJsZheKB5
Ac9nkF99i5f6qWKQHVwjvjk1mq6fzJsib2v+/12wAw6o7Os13wd0k/FBG8dSzO1oci+m/SGvdu6i
k1ohS2JD/J32zkv5ZU1SkuPBGosVanlVQXwjKOFiXF0gs3HRkjJNAwYFL68PrAiJyI2rsmVUZ5c7
ZTtLlPZ7jduXeP5JnuOOU5pZn4B80yzvl2MTB9oof5w+EFozOdAUC9ibkJKyRrnfNy6wNIvWcucK
gnWrzi5/pZPA5WnBPZFoPAdEKJsW0Td3Hazz65Rcr09rKMug4y6FRT8Zowt+3WNXG/PTS0hmorr+
48gKjpNZS1EOz/5JBXaKH/wUQHHa97xYbHQiKfJ9ZO9Q1OOImwRtkyl0AlqOjz+SZA3vOXvMeMhR
DZq5nnNxSm13G2gfgmhx0znGcUeBeGKL0lMEe0A7u912EGt9mLDhH3mLCNVNrmeFcy0ZUZ83A/Ir
NeNmy258PwW8KW4OEd6XDbi0zOTKVT7aBeEZ7HC3fZ4USzRxo+GVeGKaIV7SWv/xIcHP2yCF8rHx
5aHKdqrCkd40UBV5KLSE/8DefoMVsQtF4O3QX5mCV/D5bT86KH0jdYMHP30t1ItGXy0/fq27H5C2
pSeUFExLBmhE1dQNgWGItpS5/r6iob/jg3d1V5J6Oe+LlwczscKASfDE9B9FkgRQwK/uVNvAL32H
cxLqA994u6XexuGlHNc0Zg+vF3FI+0yAg6Sv0+zwztIYPUsFc+55FA4SlseBWo/3i2odDv/ItC4E
zS/nfO3qc0+sZzDeSPV9ugu9TTdyseAMK45LdP1NwH1xUvB8h7f4s8l3kN61D1vIJVOoYjgehzio
xexe+VlV6iZeR4xwgK26jr5PwYGMwVXVSoFSfoLIMigTebwyQXZJ8t3wu5bIYv2Jc2RzLC+anIuB
xYTX+hwqBMGzphOuepp+WJEDdbxDbJjWhQENmeB6clh3vzFfuCGPubiJ6FsyACNHzlo4F1bft+5v
bEUaig2MWjQ5ShDUf5kqvuqTYchr7FNzw0kd3WQCYUucvK3xiUF20vZmx25Yqb+LlUCWdbdaNqXd
Ry9wh3e1H64ySKJLN+y+XuEaTku1oCa83ewfTPL0UdvjtbOpeW4BqT9GlNVEaQN4Bt/6Zcs9QT45
yyqxWAzWoOcEFoMEeQ0hRqoQTc4AOBpUNEbv8gb4JAYfqWLOjysy+Wj8bEZCUSvZiiQoDtY4hBRD
7/98DlRmBWFvaC0s3OM9zmfu5tZtJyPMMR7fnDtJAGh/2Sa8jAWZJYdA7UroV5VmoXiijVfk1/yD
AlThx1iOMMdQHF6xnB7lbEqX0thHtRI580oA3Pwl+yvR4NgbhdHQdXkfd3487pH0dsKFhByirZ86
rnygzUEsimFL+TsxhiM9O1cgMfD2CdqHOFwGtGFN61CkL1tEL+8+R9bubpRhYVZMNdE9y5dEGUsg
tB1bBv1xYCY2zVXNfi6qW/sYSg/TTIGJgnC8tdh+1wE5c+yV5jsUiQLGP/6+8FtVbeO78VYXMvQb
ohlY3U1qA0Sox1fxagXCqocaFFFeRSMSVGlgrKXHrgoXUyCezQUkj2RyNkhQO/xlc8yoiN5SjbFI
j8rU4n5nUjlSQvQVqNus3PoOSkkkyNqfffgtJapgvZMAaQ0C9rZChDi2bGDC1cLn3/kOALyvsyBb
wt5omf2LPPSsmjZZTouFZlQ25mUHZTiS/u6MILbrpzdCoDJMVdvI6XI8/V3O4psO64Mw82rB3BrD
uc1/z7EOpQJH+PuQicIBCMIRqKOGwCnULnO4ixpc+oWcbOEJk3XHPxk5fcnVi9J/96R4Li6P1T8w
ArwF5bi13HbpYMjAbLaYfRjbI0LmUAQKmUrKrbgz0NKGDLen9PC/LC9BwbExb23+ZyRigwC+sakY
anRjghXMnTdQ3ZZ952+n7pqmMiL/rwFD3dF7WYE4+u5h4QdeNjL/bcKmm+G19hS5PxqRjvr3N0Qf
Xl8N1cLsrCao6VR3d+a7akemgk0kDSN3XceKKYEWAfBrnj6kQN4dUGjJ0RR0aJMm1+Z/bAhuJtJh
OaiCPeCdBFFYRPyQB4I6qWtikYRWYcMvO7r/ZK4352duas9+Ptt4zE0CBVCtk9eSrT9GS6EksOXw
CdBB69khpYwCp8KqkN8NMVZTctuBkd0k8x/5yNKJt6oDYZMEKtUhOT7LyHi11qNKn4vnvHMb79tM
dW7QE8vSzqq4M4uj+PyVbwdZs78wK2YfkB35l+iozYJelQ4XWfm82ARBccWysKBpN1paTYQxuTfm
6tpnCHyQvPd/diy96ZOrSIxzQxtCNkLT1ZN6/4MQJjl/uwy4naPt8+lzsEXFZDHIsdZAzbY4YXN3
RE/7YqMPgY8yGRCLM67MGUKkozDM+Ugtr3AD8gUyoa7WcSMbW0c4HnSIfTzfcwu+yym0ELAjJ/hu
JJVCx2JTXkbm7gd3wJYss/x9KATXGotsQCYnyjvLN7ZjMwrwCcrNsaLTBrJQjHLBH4P/uWcB7dS4
VFKwesIC3pYOKWMqO4DgDvLIqZ5bU/2YDctc4UVk15TzPkjkp+A44DbIYYtlpgQFzyOys4Ou0Y/L
LUU5rqYayDTShZLm4ehkS0eRMl/HYxGR75l1Or5+fq3lmHQXn2J7jsMVbpl5h9fBH6+0njvUNaDy
fUS4aKktTympH5cnmwrMPIPUgikTIRSzEtWusotgPkBlU3TbezOUKg84L8SJB4QDFl8fnL+cDnLX
xTcEwtzMHm9FGSsA43Dpks69GZJZNyoHftiqGdKsEaIsvKpZjUcEul1M4WLoSEvh20QEoxwSPMCi
DtxcmfYLF9u6ihsE/zl28FeDD5Wq7w+/wYu8fXaTrkcVkK3iLkKFQNOX8YXgyzjlkU7b/tR2KmY9
lJPDPLNkHLdWM305LETKJ6xwwtGqu+EZzoscHXC5jtiS9wCtqionqTz0iI/YFHd9xbMjmhJmixAH
8TPVEjSG49wcGlBQBPf0Aqf9YF5kXewO8IUKJJWwXUrIW46zoRErRkBb0wsGEMgykO0yxNa8u0VN
hI5vJJ4ZkBiO/+ixxieSnQqOyid7o5cif3zp/3dbeoX7q3bqKJbujAr6avvq2u6XUGEIlLTlfJuE
uQFE/5UR+BBDMrKWh9Yv5TmFU8pa+LYEK3XAI8g/8IF8N57bw1AMPkw8dHOoIj5kemROk2ImCibV
tSXkHc+/2Y5PjojkQ41OpSylUn9zT5dqNAut0a7n+JcbhWeRVYqs+7+PustUY3u0K6qPTPAlUua2
80q3fvF6EzlUdTX2G47W2TJa9q8/Y61XQd0lxW0dKNTwJSuU5D9h8VCkKwSgifWf1va7BrFzXzOK
IPxoy78+xJbOzePCETjcCSloPVOkQZTsswwtoyMiL4uKqd98nNWA0SYe5+QBHRpM0zWu7Qulbmjl
up1j56led2SWMwxQn0IO7RpWahzBxxra8ecSKvyL9uFHxY9VkccmiPUdCLybJBv8IATPXllcWLuM
USGRUFtWas+efDFG5pDN088CgFRiMSfqHYSTZ5NfY117Vd9133fArFNit98wDrOup4o8SBwPFVVN
3B1DoCqSx7Sob7SbvhQtlBmS1q6Nq/UmKZZtVJ5bJaEZJm3RTI0eWmCuBszLgYP74C6uk3jNnp5T
njg88HnyueRD/eUUKVgWyFJ8GCIM5qVXK5eNkMAXm0Xrt6LGcVbBzoSeumD58ELu8tvAFGPI9GAe
5wSZbiiBtzezv/3dQe0c9wzYKtK9tJOev5zMsNcfIeQ46xlOgyryUJRNOVbrMKInEjJ7u0eOrAfW
Acht4+CLCictMtBsJQb38KPGS+oc9JEyjSgveDlAh+M1T/+xjhBXOMnhnTyPBqmrsOiCZj7+nGIo
1R6lJnz4e1c6IQE8wwL2SDqF0i/+mrABluWUyUGdDdm+hVLaLx+O7c61IA9bL1Ty8PlqBjo3myCl
/LR6s8bWOCnJU6tvkInJ4hLkQb/EU0QHWDdyHoilyLR3t879BS3Ns6cYKJL9av5vns2yCjz2qbju
MrDcnVKuN6pralHrxXEyxeRGtKkDjHYA41X/jHuZT2Rw0NVeixA5mTpBXUF32X1MlktpAqEnpWm6
r4Ut735yqnSMAnUvSMMrLBTdElnmajM+UG6JPMyI0nz8Oezz8VUYfpUeCTR/EwIqTIM+6b4G/duz
rs+UfJLMyad1UAtf/ZoL5cms1kKOPAOyy8XnHqsjV8f+mUeGHrx3nzGJJd2/b1YUBhlcBX/dAHQH
5hrw8lMKtsahK2YPxnwxhOFGWWr0C6Rzlh+zTPJ5dIAAyGetbxXofxF47UDV7yLZTgnx/rKE7QPA
QvVM9sV+YH4k3NBC0Agw56yq8kjIedVXQ9O2r9FIJKg97AZAqdBL0S9SoluNmHI4jFPUKcpqJ8Kn
xozPSkcX+OBt1liM7XmVv+Dx+lRSLshyRDKyh3sm2IA3Ehw4h8FVDPl+pkGMyLH1jGQbEiTqRP5a
b3XvM//Qj6qW3FXf2s0YDaVVinWTMvw0chZE89KamvnOyb4H0jE7AkgJ2IuVE2Ggeylz61j7W0Hy
eI+yoTdO4jQv0vEBaqI59cVSWmIfXDBcccrbJcE/H+4PHx9qVtYL/dzjKxhDthxg5SczVWMBxYh8
9iOAs+ACpLZBBOvx5mYeqYDOfMDCrc1PqAsYwQHZ+6Xhp6/bmBKBNrVzbJ1S1pFuVj4Qcgxd3grG
wP7T/0RRL9jDnlkt6NbFqt8LCdi4ezkH2At2UU7yNH2UVX33Z0rvEMngiOef2dPzz64mPQzB0+ti
L7YxplR3lB8fGtmnMbVP2mu+dIzXPckTnEaehu35aHWJ7n5x23VEs6dphsLAyI/yDMqBunOS22wu
ipMVRCkyeTxS7Do73AeU0nqpy09o2FeZqNWX3Qptam4gp8CABDlr7ApI8mHytqIWH0BoPX0zxN3d
33vItTH69558ONba27yvDw/gm3PR6eghwpOHPJuzxM8v2exTa6XnSMoRkA4yGKIPkZQbjTXfhln/
FGzDDrKD2B1i7ZM3YazuAUwCpSckhJKaho2O2g3cGimsbhXb372STQrSzKe9cDd5LUXYsHsYfZ4b
FP3UK9Ub9eHWSWCK7UawNVi+a6uf/lnMmvoLU4yNPuG2ZEcnTf+/peMbBbdWYd4aP8FaxnyJb/UY
9bBk6ANnV6/8pnDwaU1thNPfaJdXzjp4LlaAJSr8oobxDOaPy4vjfNF7AC1RzHgRfELaKWS+Escw
LV+vpd3fOaoL9HkssyVzbf888YeRgFgJAczqDW3zB82/+f4LkiD9wMgc/Ws9ijyBGVpln9ZhPQBE
hxM037ytty0SRW6naWzjLd5YvtDJZN2vYE9v87fAUxEoMC6QEorLX/hW6KteXlK+MVAPD1QbPuF9
HRRBNBb0uQ7MXlDwYmjDIbCtPAnlHPfRJTWdV0R5RaXNo1As1WyIYgRJqZTqRnrhennB5uzLv/39
aHyxvCbABobYbdflf0F5uNNPyccepiYkw+qRQEa1zEhCY5/9gn9ASa4T8VGPw2nEj5JXTFEIl+62
1uo8r2xaukveF4qj0weF+k2C62SNiIIj5MSXcKkaIMUin+aEXL3EKiwZMQFIT/QmAIdU5YXebS+n
JLQ99SBhSIZp8F2XrBkRUTlwnBV30DzTJl3v47q7vp9fR0Z9W8fK5jmR3LGE0dkxxe7E/zKsBmlQ
L0n4/8ppVwmFbkLqUpOXCas/WsD8H7LMtwhmu4vchMd0K/Bbmkl9SrQLf2x6nJn9tp3/Wmic1gEY
x1srGSY3DqlgLR0G/gEKran6YGiey4VHsH5Fuo6q0PMg7ixHWr/aMFzt+uPMS31b9HXhH+HtF69M
0sxbEv+fbMMcZ4U5g/AjOMm2wHzN/fvP6189GlgBzPPo+XlZRWdPk3pWd+kKrK+Lb7elwyxgown7
SYb1QRREf+SGc1XUUpYkPg1t5gm+Wdu5GtYwtT9w2LfoS2EMjeqrFeJS7bncvh45c+BorcblIAB3
RdZDkuAmccnUsFXTeJneFCRtQ6vYkv7LV8C8MlbQ3zRQtOMfmLkI8e3CbqhuOE15On2mvVoYt+h1
qAejhKYdeNPPzFKv8//mjGTdFrm6AutCPYWEzLp1zHg1e51tNgb9IBjEAFikdfM5DmovNhDRHkuE
YONnZcGt9YbkImsPUPDVgm2N7Qlp1dNyzp50Bqr/5+KWuUP5oMzPWLvpMdig1TzcxsfgbDFT/uPa
qWFwEX81/jLnO7UGpVJDSnvVZP8IQtfLbKVBXWnmbUES8TykBudihcs17088/jG9kZBldIVB8klR
8SobvUXYCzzA249gJ54sYRM6LNZuOYj6Yjq5u8aY8QrY9pyW2Kz7wRH4IWWGBSKNfvaMCunjF41L
BOFNkA2e+ClOkeG5Vwp+9SFALj8GydgW+QGKXG2OALhzCsCiOAd7+46XVJF2foLq/EnCmwGBt91B
MK3/BZV37vwU+PyLFQ/IYwTVUqAN3Js/r3Pan2mdBpywu3G7u+MCrRmwOqYwrtsrwN88TovoxMqb
74gYPULFTvPUZDZhT9/ppBe7UPm7DTXpf3alFQtgyTcJPtxmeZs7VgZOVNtZgzmU1RS2izIF5fgc
iBj5t0bvWiSXLPaz+3REnOPvNVN3MHC1RkryZ5308ERR+A6MR4Sc92uTg5C14IIy+L+OM2ett4Il
worWVAEQLQ+aeaUsDGJZ5p/9exqDGgqlle8zJ0YoQAU+ySxk8NxoO9wNrj10t2j60z2Ye9GroAAg
Jmzwifl5b86PuNAkzVSptxT1sI0ERCsBLVKczW2POKtml3iIhXO3C1hk/xz2pNLcG8pc2UO2rQmC
yqVV+cIPnbR+gAjoBbiWzCqlleppCaLPSpmuRbtAXNSWEahtq+CupHopCoVbnZEdjjzws9TApxxy
ehWWlBB8i5s66IN/MhOjatLo78UhAYTZ+mDrMrJHKUCKArUX6SIk0PgaFFFF1A9WL3Kz2C17KgAQ
MrmXzPsBoNrNZwUZ8npqX2txzAJAfYtjQeKfgolqU96LASVCRhUuKdIaJG9SDX+MZSBMdIa/zWEy
giFVZsQOJaYGEgyye2kMJx+HifNkXc8VDZEXf150iP0W7ppRrQ1xY1LjPkEmXUwBraGeSjafuPPX
X24u3U78mAAy2l1f4ZmMvt1Px5sk7YW/U/qFun59XuNH1TlBvqBl1PUgjYQocXy0Rr4Kg4V4yiMq
LaRb3ohhhTIxElHwAPbQRY4MS/l0ZbeMtNrqRXIrbuYgopjlp871KgBmlQzr5w01Q4upx0HrUU7h
xTJiX29lMdrRES/kUQeWRhUDTVw4ZMxjdBclJAKXt0g+MmN/oVHMsk3hdcDbNJueVCN2sKYgKkbR
aAWB6c9WD0vsg8VY/6LThRbS1HUXG8fM2wojyBba7r5uOXN83xP0P5YG57szSlcZSh24UrAHXVLD
gHZKMnQN3ZE00K3wBMKCmsSiyHOGH9g01dFq5rmthPQp/vxr0qbPjJE242ADrmBc/yr4qmgHR7Oq
kU4wv1KvYToxRshqGWYqYBU6iumPAHAPSvsaAAvqAPPp+cR+uKMknZKbJ3yn2SbjnD18pg4TkGzw
TmcpI+8mYdntsgWkoEup/6uWMfm98t4yjB2zLKq7OIe8WovGgzEZTO4S/TQs7V7HrAgUKvS8UlsK
jiJA4yPFsyOReR+BnsOrihv9kMyFAh1C+5iAIvYKhFDZYO36xfZBPHEDV3hklMDPbwSBjn1W2vsA
ygt0fl+/RUWcxaycoNaAyo/JuuwPleIngr5l34LETP3SKeqOYCLVlvbtL0K+qSK40czlyflxC0Ws
y07pGYEpiOat8UsXyHuhrtoQnEXSmO9MnSCPJ/mzwUdUwgsLH0acZC20fLe5E56nM925NhqQDwpM
fxcEOWLHg3DJMDd2Yfd9461bIDohKY3OWKjde7ktPngedQf4sIQBMdOBLKV4FFD3n8EhQxq76z8B
ufuUo0JkUJXYf/Tb+eWwrE3QcZqPkUDO8UU22aXoxqVhgePEy5hqu7FAZu45+BTmxJzs5ofYUGV6
YkFovzC7VUTvc+noi4WaU1sujDoRh29OVVpJoo0eynz4AG09D2g93UhYAmgCctKGm7TcKYRI752L
4vmFSfkT5aPBKBQjqy7TobvImnBOUV0wE7bNG3yYYuEW6I5KxNsnoH63qL+dQj6zYloNwYWojSw7
Lb1BIKGcSd4ggGySbgoRxAoKPwvUZooMTNqmBHpxEEWoOmOLZtSACwNMbfDCubdWM4/du0bRdbjV
fdkFeftdKAxtHm05vt6ZUPH0v+dqSWskmmydB12Bzg4B+hxoH4GvSPO0dJgBqrHmwV69Xjfufv0D
cp+klrBnBBkVgXh7uX0CdkRqfP+yq+OTswpZFicE3A3mZJD5gYoZ6FyPzJCupehOhR7MPO1kRkzm
BljVouX0Dm+l2c9Z9/1S4fVqt0++dyW9U1Q3c1zY4zsCoH4zN8/R958rJJOLxi+MLFcBcN5xPfcJ
QzIrt3AivlFVRYUS5F9W9KzDSwbbd7q4IFgkdR5qnBFFHVZMIxcEUZi1BfcZcIGg63Nrk9YAGqpc
0DZJ6uIcW0SrnhQZrd6UwQgMy8Ghh3hohc4XXp7Iy8bbP92TwPmQoP3bH9s8iR/YBV5aE/5FtTjB
BW+geWu8C6DcG+TBpuPLjuLVx6yaSHg1J+pj4t5fBnVoXp3xaMNoR3uBnDjuyi0gbQ6WogSiLfD8
DWM4IZUKnNaj5fi3VH+yLegXDYjqgnJdATURp9v5AmeOIF+LHVQVNp65BDSosvJRWbw3MZqGoToq
lIttz/hPTMm6Q7t2Zu5fiIaKHQ1IyZ6/3upEMKVfkZgUzPoZD8ehdJDUJNI1gKbjwznBuFQrMetX
djLJKm8y+J71QAc5L5k6t0bJZ0eNdUAFyScA7xlD1VMtmu4G2W19pXbILxYly+Yc51pIxwx65leG
ib7hi6h9Ooion9R5IVTTi/tEbkH1gakxs9VpIb10IEjYn0kZkIA0M3EJYFG/xIedixrPo2vVU2Ve
pysK3h3rbV8chKnppvAsg+GPu+ejfsWyQDLP1IR1FuToY6zszAP9aFIMSr00xs/Z/dogkp3YtmqV
Cq9sjTy06eAGhFQk4gGchhkl3cKeZ4Z0ttnYCG06JT6og2/D5hMb2aq9grX/DyA6QoZPckAtFWVT
030qvDJ8nRIvDPHWVe3JMUrZqlzjBwbnOdy6+OKIlQGy+YOx1tbmTzwtFd+Xyu42RAASUXx+j5ST
ASVwFXsoG0QdwZ27w4t5XFb0X0kHbaTYrewtk51Iu2RGJ+ZnpE6DpeLST+pg2Ix+ET+DU7R9LcNc
DB0b5pIq4h0NGqb0/ZBCxQshoDIwRD0DNLmWmR7VmWNWwizACtuzV1z3vXIHf8VEoMwfA9YHWmf/
Hqp24Maka1MD4OSPlyU5ryMlVlMmUd3gBxCyGe/DdyYCDooz/gFmzcDQocDgjoimLzHr6xynsk4Q
q8Wmj2tHnZa+9d10u8uwNVrHSgRm5uZornry46mmV+yAPm7IZgtnUaprpiBDLs5SdOF/iMkmqHIE
ev0UfaIqeVmVSxkr400TcwVRaJQTV0q7siIyrjdrQk5c/Zvwrm+bMnIKHg2FP20lYgMTiryXPMw2
6Gfsa+0jaP7nSe+lVbQcT174B8uMvGhYEq0q/+RWwDXYQf/jjkKUke73CcXTdoMtvH9TJ080CNBK
bH2X58T4VQuBM2GjKZ0FURrEMJXWn34JhxMbyqgU+ygsT3LFZ7fbvfz7Ai9iKJWTPnFqDyXxLYth
zKvmgYTbqFJjwCwrHBMcA6jg0zME+f3CQTMQhQEtiBLEwVf1JTAF5AMMChew9+7vHEboZlDnXAga
NSvAtUL5+6E1uKd+mU8EUPVpyWOQFGFjUkC6tq5vJW2o4yYeE6lDYCY3H/q0TahUuuFA0Sxm9lKe
BoP7sPxj9Kupfwd+fMl22ww2sMYXsTNnkQV1in123ndFVgqMXmUM7a6KBgAuGuNjXdwuk17MmtUx
whzSYQ2aEKXlzmQGZsULt7IVABEhPNBOxNiu1j2GU/fK58XrBRuDYR3b3sdjO7ulwzqiMUDVn2tb
hRzJcCmKHNEHBCf1kVE4saYL6d5W1RbEAQREsQWuSfCgnSNCgCGL/zyaCpi2FmmkSYKklSfL4sAN
iYjESeLtx/P03jBV3G93+LghGSAhMof5gZuQ9jN16Ay3aCR9/7BonORTqhBzsVQLVhCCQu4hzaUD
r3q3HmFN5IXXtiIoNUfd9RBiYeRgTsvFIYTCsgbLRF1+PN5y0a8TtFLZNbuqpVIy4sqgtgZhTwcP
CKSkgg7IyjQsHNSsJ3Al+tASJXntXLeGYm34y2Oj3+NtWNE7uZs1LO/9UxX1nJsU44VUJNoSkEhH
LSvWsR+KRU5SikVsnMJ/5Bk82W8NHWRp0NMHxo4UOOBJoj+1WNh05zWlOlCc1sGwC/IdBrQLxPD+
ozZL5HRjIBsArcFFy2f96A8QsamSUWtLlfsmEovfLIhuTYksR0KzzasqvqmvDaj1zDo18kSvz7on
SRhVGKcC0nBlfIr1TRscQDvQk+iWbdXgRRD7KBNFHaeT1ce6Ba3sUIh8pUjPcffPvSq0rjxODhsK
51X9caUVVQ7VXcKRpUQCIs7uJWVTuoWivBLjsDGbOl3wepQbbfnwueoPqscuhiGV4XTDZI2BDKzy
BEW+iIPcF1nORKdo1zjeUhwAMQ5Iu2SRQnAwLuUTeGrC/5mI1sPNp/JfVQh8ssXyxNFzMvSuHmpT
ZnfqYoUxO2Mw6US569hQqvUzrArUPEc24QsK9PaQlk4OhUF85dXr5U39vKi8CeWxhydwAloAK/xm
zIgO1I77vwVu6IHLXanpoYFeCC1Z9lW0dFrudizorYY2NZl5OV+fznPetlw5bbqksCTW5CO/zfHX
cmeZ088/uGggmrY/EZAL9T4waxO0ggAhAGtBZeLkDI969EJhFcYnKWph20Q6Kay9rzJ4Q7q1Ye6S
Je1rtqNp6E3x6aHd+rVYT47l5hZ7BG3+81eKS7ivB4EbphMKeJX7Y72T6IE00eL+qteRg3GnnJXH
uJpseirmG+KjG0f8pwDTTVtBNZb2pXAvRSxwMI/jn5u1TYNYMZRbz6JxwrT72YV+Gi7e/UUYEPD/
KEEdaHhlXexDtxcGLvcrbaEG/rQMZzkwf7bUqtAheDRmIsATSpSK/R1SflD1fb7/1HYDEVNG8sD2
EpyUvpZbY/6GWGQIqJzhu2/70EojZUrWDPZKWTVI1RlWsyWo8JvvZ0IBA5QMMLa0JccHGrdtrKIo
c/+ApN1V//EJQ6PWax0mzmG03fceMqhqugu6PdiAwclAd3sB9kgt+ClUb5ROcrNjzQ/bcfm00stx
2EaZG2mRA9ZqWeArDyqEfHSAZlnSHCx25XYRNA1BGdfQAuiy/D2K8eIVsTtYT3OFQliKq8G1RHwy
51B1qjExAg8w65GFULsdYHL4XoNwHnh9p/VyQPxq+NOsO+h70wxhyvzl+btb/OybmmvSVOrD5gNZ
8unWXxQGwB/ocNLsHwMMhskLW9tAlF6p+bQJ7Sc9oSa6DxsSIKYP8bdvxDc6GzwQ5aPtRbrx4y+N
kp4JE0rcmRevSG/Pi0kNt8PvsPOgHl70qTVfIkSYehHnEz+B3DBju6yzOsrabU9EGuamWx+2/txw
TU/SLddW/UKhAXmWz8z2+nLWxXrBTymslK2wGEYY+vHGNI0NnZ8XRKig/w6Gpj5GKGgWXQGGSp6P
hjcY8T/+nwTI2MkrjJD3PNnBpce2uUEhcFmt2zsNEkiEZkE1m7217i4q9R5cSB+4byfZZpZTJS5Z
+X/ZYOayrOi2Jl9CvNd8es0qXWi7YBtMcbdiGk8u0tJMJbu8Gle4Bn2rqUjQvvmdMUU74R+j5aGo
fMcSZChavY6RVYRavN5IkE9FN/KKXHDuh+3OxtOo2yHCF2Kr7XHBmmFUs3vjlpdr8U9k+p+Dsegr
eZXK5enj2amNYp6x6gnGLnRhbhiiYEWvEv+/6fxphz8lcJtrVWCrmRvmay4PwWJU6MUCpY5RyKf+
4Ggqc7/JYXd9xTS0kF2fNT+c0URwDfpLy4K0R0uW/nj7TLEsBF4LJcwof/0+UtP+KtGf63txeUrX
I+OK4bFYFN3TpP2UPeV8q7YaL6fAvbacgX6GWp1KJ0HTF7NWbRWyHRKJ/H6nt/x/Qn8D5bQsXHc3
nVkr9ch8UDsfHD7Z9IOGm4jKZfKGHkWbNBGa6L0wPkcX0NSDtPcRDeYEZ5RuaYhjRpIXyEQoLlOA
uSge4mgsVaI1Lg6sSv+uOpe448jNPJerLN/oCUDSFkuQFoC5EuzIxd7t++Bvpt+2Rl7jnOiEOSDD
nKErbeUaNVDkZ3TzY7OOBXMg73PWGepsD6Y2pbrLsOLP3D59zqZSfvpv1d5kZzohe5RtmQMLHiQe
hk+nRbFfbJF/JYuqqMPGRBLIA4UdwFJzgawnWC8+fo/7hMjpasuQMq9t9NC1XAVxxJBulXda4WwW
fgMJXcFgGaHRPmiEogz7P39ANfik9CaIdiYbd3bx+4iFUHSWtJw9TixxVWjHhKRTjxHCwL5VAZkb
UdE1IDe6Hg23mudCRsHuHnS0K0OOk9DCF+fz5uM/i6eakqWLtrH8koD5bi7wmeeUuFQVPTj9L/Qv
vhwxeDfuwul1Fy0AmeYHYCY6SeW9MikvVq0sbdDp02pZhJvbwM9ytpzk9jVGRwK1314OW/BnSpL6
a8knOlL6TsQJLt3hm8qSRZv4QMAgATb+l5oR4ECtbWv+rGoe4Isx0NFBE9LUKqaNkjuwKn0Nzj2U
4YAFB338nwzftikhUtKczrknARy2ueK4oFk/GBCgqsHKohfg2ImWZqPpEVmY24CSeAG8g810+Bsb
PEH9MeI5W7nWjYYDOOzFzFz/lo7H05CXpTxSO9QsYunlTrovXJYfieWJo6m3UIy5Md5q+yiFkETF
1MsjZZ2L8XLaemujiBLGiMbtjwVec6/FYqTxRwepKpM71J0oSwP5biks6den6xSahrqcauynZ0wn
qK3+tKi2cMB/tJxGIAj+6JvClvI5V33loTTNJ2RgW2fS/jCHvekeV5/29c7wdiyofBmqJu5IZe2y
bFS/qn4wHbT9TzQT2eMxD6gcq21lQ8Pr6O16NiHJ6xlD830Qu4kw4HZ0g0Eg3sZ0Z2tchxq59T5G
ts6ntqkzxHL/F3UbsIlX+d9IpQFdeaKaQ4e3s5lTkYneO5HtBIwbv3nETGKE5SRzqxZ5JzXmhKn+
TD3KGUrbU/ZVUmVFzfmTLljW0EzwAloDv7HJKt+fJXDyLg1k5pab4VaVh8BHvEacmrtNxUXVZTzx
XDDK/ndDrRLUiBamCmW5x3++Z9LnzhGBDCyhPPuV+3bquG6gVGktG4u3F0OzhrnRAZHmg+hSgvmd
D/OFGAlNndN1R9Av1Bvdqw2txhSDB1XwSE2JLD/7mbY/yFlGZRj7EDoOv33ATHtS1fwnBd+BtZVc
A+yfVGSJyr7wxpqzR0BTU+qpnYm7CDNT4IqSPLaXIjznnsk5hvdLWC3pblfgmPdZ7enNQXS+rtzb
ync4gJ1jvp9Nhb2UqTL3vYq3KzkXVkWclgK/OO80fJuVxjPfgeg6UY2vIJgVF+4RbUnIhlQ7RFzK
XcpkFnRCihNx8+luZUiqGhTIrdf5HQint+X4dNOQ/U+A+vJ/v3/rk80nbtONah1sZhIyFf1xpcmo
UCEVGlupxqIp7S/Dj/TBpoAJui8Wh2mpr/9irOVBOyct8MfWzudDIyEWNokqO8Q7hLo+9mWnBuh/
HVu6JiJxyXk1m5jDUy3dn2d+3sVKh8+1lzOeo9LtNMJXFLAPylwuKZ1zLPD2KF8JqmzR99vL2NUP
lGRstThbiQFor+dY+4e/N3OixGKF3m7pTST6PddWmIez/oXcUhHDaZoOr8noKmIn2epnBquRgbCK
TT+39MCMdF1uBgShwiWlZXZgTD72Ayxaq2MaAHnek1391OOlxPG5V/O3/xSrVilNBb3En1jJLrH2
zpkPRBMO6wS0CsE90HB645eMQpU1fMzAUvFc4+ErUGZyNJxUXbpQg3le1NTQ7T1XDdufATWW+3qc
dj12A+ZleNOcoZx74kacLI++67x5UaF8Xd/X5iZ18WX7Co+K0PBJUqihC/ye80VKQWI/3QdPuHwJ
2Fz/kzH/SM/xXMbRqmOMTkjIoWRhvuWfIuRtBbyzauezMxKPopAFm4ThbY+9KDTEa0HdhccQgzZg
qNqm9m1NBpGXj0QN5+jzxjI9deLC5ToaEjNWLYIly3YduIhkQu07rdjfcCMSUsbrSK34wOp/+JM2
eKIbHzY054xUrrEnJSTKzFVen/sUacjpbYLFgtsJiOVmzf05BAdQBv8qkc9xdye94qzk9rTlnaTk
saSiJDcogRbQImG4wW2Li63dYzCyGtx2HLL0FgZV6GJGqRJRcYwKSGvTbviVW5GlJR+v2sSEt+Fu
IXdlBE/J3Z2e9e8+yIk+I+ssA4OR26xR+cPcXvcapf4jbrMpAj7NXv7b2Dup5ItLMkKKIvH3vqIq
ll3hMCWn8frWEY30PDPHfvl78s5MoQSDHRRGptAAwNWPXPI9UevGx6L7ITDiVfAinQVaH4/Tv6nQ
ewsWZ17ywRHvRboCisqEFwq7kslRTc78eZVCv/xCO/IWIGZ8sduVSiKY0W/+RswgnN4wRryN/oP+
MYbG4CV2PGzW+emtZlyD0z7OlpP5qTAeKOGw6rIJwdLdFdjBuypbtHrJAEwe08LKf369gml3/Jur
1RqSLGgGNEEmp55pYuIDIUDYASx7xbjoLcToB9TaE/gGOhZzXMj+A/HbfpzkCMxjsDsOa8eOTLU8
WwszBLP5UtsLjL2F8EqN6ahctahtHizksAOLz4byf/MTNNIUkyZVLPsLt/tfzOsF8o5PMhAu2UBh
1HZG9PAban64kXP+vtU21m6ObUPTon/bUqkB2sF3pB0TOEuL66u+gVaz55MbMQexMikYQGOpiclY
LfrGhEMtJfQG4RBqzpXvf2A/qjmmdAe8PNt7gHUU4e9rlirb/c+cswWEdSHX311cDiQ6mYy9GFkw
A71DMASwh5rypcRgibrt2W7wYOHWU/LhmOuQgmpDjmBuzjHYMRCWVXlczStSCZvCMWd+AkE2T79F
PgUx43ysAZGj2HvwLVHLr+ZIemS+UovMBBlJF8fo86vi76miXlDKbVyJD1v87sJFfAaKZ1RkNDnr
7VzDmx4WNlXIm/wZoqoJd4wO90ApoOBd8ZpNAoGICS7I5qtncJ9ZM2pH60JOAg+boeSaiu73YW9S
gJVDzgBanFrvLNITQ13mFYiRrRcdOVpk2yGP7oSHogS1vPq97f72ASkUZPJxDpzgx7KbOf3bSexv
Zmq1E7y5CoyTKg4lGc274/cI4hPJ4hh3zZ4aUSzBsDVGvUDRkepf4URSlC4JC5zRTeI6gPfMXcRs
Krv0RZxA0D5CCA4+00EpdudCmZqmUhPg3gNxDh1Si1B/wHmxWi95STyr+K9OEA4f6xXETLM56clt
6iEQ6ts+4OPgu+psclZd65GQQfouNCMpoNP7sFvAgsEbGB15QWMGefpHrWy0A7AKgE4/9wqwRgLs
cAOoKPhRSq8GzqnacU15/jNTOwxmGue68R4mT5KsdHJOQZpx8Zsm/fdTZWpe1coq7+oPdMXvPMFY
C5oNLh1PxOy9ZzvgXmG9pOFEjQBZDV9EgO5nU4vhLXhACfOVDzmKvyFhK1u+MnUppmW420KgdiGr
fmLqfh7qNlORclLOK0hCArPuWqfzisgF+KSZxU79caRZaDT7FnbkzIIS+5gHIngNNOIz7yUdXSUV
8uqR7iWIc530Ihz/sLuaXSOQW1pt0eblt9npjzFh9zfxfa+0LqCu0ANKXgYQhqZj+D8UIcj46XvF
WtZ5/aECxGonFfYC7DDKCxnbT6pigO1SQJc12lPwjH45fHwflEU93pQLEq0hax8QSgqiSXUsSMIU
PxKQPvPnFiytYLfgpLViHL/BD7WfyB9he9AxYnaSvpDGHinDpcanF55XEu26fW/g2SiWTKzTghCO
hZk05u/TYalp23Z44lL0JDAL8euEG99HieRFno811C5vP56qFOgIlHu4lFyEHp7vF3z7aQoJeJ2N
ZQbJROiV4mNtrA5LyZgj/jwOdWl5L72dhq/YUaqFl3T2kq92XwCAnnH7aZVg8R0juIyJIDc0itTB
bx/TiezUeZ3SnXJE/9PFfD2/JfUu71maRmM5onL9daNH3iobaZ90EdV/+3qsAw/VRrH6qyvpeNov
iHUE61uMOKiC5/wXVg4K+zMlb9xGSu6/ldJnydkRFLT5Ga0IOvwuqVaiGCX4ui3z47e/D3bZtTeu
R/VfrL8bEEAHm7LOZJM6el46Y2gcz8H0R8RrbKx+gv9KYsGBS3BOCugedq8n0AyAfTt9hp2y4nXF
Zbu5PPrZq1Ibui6CaHbJeNoISTBygfaBMEo175+M3PMbYRRuO1BRQbv5/2Bq3hHMUVxR8Kce9DyK
Ljnyovf883PWUtojt+KyACwwT6F7sqUDAiQ3hnXzY7tceOqTZ65CF0rv3cz3qqBqpYElTNnjNJcd
xrxMj34hGx3kWVfuIq7uR+A1MJh8X2cbqDFk6pwJW7q5r5nhGPGec2j+1mLA8YETYLJczSZX/zez
rGRqIJD/wt6ZWaphQ4oGJeS4urI0DM4VBIHDMc742mXl5MF8fOL2xhW3aakFEhFeCAedn/9HH382
NvO+1HPC05C1J72I1c4EvuwwXZEtbq2wB4s84U9hywauZsDQORHMVwUBl5EhL1hKXiVVDlh6Z0p9
V7TCfq1dDYrmUiwwUR4sUPOlDUQ7VDit5Vz8Wr06AOldbeKpiXhSnllB/+muUTOBvKt2YdpZ7+HP
+NOwFQfRiIqzbO4kbCCsRzTFoD/q0SJAt05gyoGA5KwtIIx/OE4aw2I6DRh95cmM7azhuNmSsTS3
YXit77g3D9HnkAxkbfAC1C6QkVZHacF3/dXjqmug0nw02FvRuBHLX8tBWZcVt0Q6u+9LXbHmNZe3
3gw+BSlGnU/W8/ulBPZl1enL7Awo83mYEmX8P9lk3yPf6u088GxL0tjRTGprFAJp/TKLEx9aArnb
fvWm3VQMlTkOhVZQ0Q50pnOrVyq4KsVwL4wuypnDx7Xod9zpWfvXQZJ4xVEjc16ZqlB8PyfiHGfs
7sRBnfaxGgmZobYuLgIV8ug6UzxTqlf4E7qMFq6DYA8pTtScYiRZeE0/3iGyEof7Xj6nGNls8sGp
2LYQ2AXkdvpsK7BIFgGrPchc/C6PuFvuvz3le5dCxOHBL09nvhKoGwl42W+SAW+S/r0ZhtyWzlGQ
KFjHOK+A28PuVknLMefo4W3mYrCMR1rECdVtvoMuXVqGBTyfkeX/hau+i3UGKOYU06+boLi59e5z
55INIz1I0fGMiaNOciq0B8M5QGQ2B3sqy+jfysss8v5QBbt2lvk+fGH5QTQOgdnaCNdddfke8kNb
/K8DRe6RsrOuwGC4VxWU41K4PeacQlvsw4R91shjy/iwT6dAI8TWh1gfiNET1WB7wKvaCr5l0wSt
/Wa92C/dHNS22nS26C7/z928g4yNMUhBG/aqZBJGoQi/zI4h4en/gECKmQvbKXxJ3yub62vNeg2a
Z7q5yZSRl6Qedfb63Hi+G6PD047Z4CqAYztwTNs8CI1TqnAbwXBdK5GAcNGkGl9mgMZBeuhQRJgE
RLFEshYTb4JqFQ5jTQJoH4upzQFbJ+ebO6tR5MbNwf9gpv24xSZK9SL0h4lKJvtvZ7JIiXuycj8N
vPkZnuKLEqHueEo2cLne1PDYXhENuuUUQ6AVR023F3pReej+uoS5v3uELcgmXIVDWOQdS76vMXv1
QgQE2ApGCT52jxduuAn8WC4VBB1qkEp34WvMjaqaAyRKnLwmyvqyRsXTdFG98qdlIKtPfgchXAd8
ZFCykTwt/Gl8o1113Pj+MFsaHttYYPduNEOR9IrX+tb15brVOnpyVbni2kVSkkl4DkzWQreUXLSo
jUJP87vuoRfYU4I2WSLwH4Y1ftZakwiYbM+f2nEqtbKb1yURibd/kM3+qurXD/4W9kpKrIMtAoWL
HOXjfpiTCV1BnVhOF7homYRx2ELQ+iI4M+L/2KGEoMraTypPQ8sKIJ3eJIpJTg+8rVvW4sxPOs9x
na9ZssWtpV8O6qPr+pBIpLLlvrC0Kcx5FUhOA2pRsJhhgS2MKDZu4q+buF3NjV+bis5Dc39F8Lgl
tVKffrTeTT0AY2mDKwbXrhn79KVB8lQsEsQWAgVPzKjgxIW2Cf1IaUNsS6I4NCP0PP6874ftsUGF
wBnSLSCI/86gzmwf/HpmtNN6z2ieM/5uBZyZ0okBnIS4wMnr7breXWGT+SIVLLO17gbSlHn7fV8l
k0cZ+5QkODdPpPAVql2ZykMHveTAn7+jbpbWm/M814VSQ4UxOZvIiB0rI7NUa82piw1gK3wDP+JS
HwOwpNs9BGl+MAgpJb8fdvd4YqTM7TzRHK/X47hkB6+EHlJQM/REITeuIFJKmnMAGzUeAYNNQ/wO
qe+JtZ739GRt2Kv2Lt4SM7aMI9VhqbM41EM+pvCz9nnRPaLCTYX3bR5pNyIQ+ZL1ixHshVlos1v7
qGn1olfS2O6YsAVUY2u1fNIOLp88/BkaIS1X2jVDSQGn/W9uoYgtOnUCwLqdQrk7w9/BZwlr7Zdf
pFXtxB0M2ofGVtXJILuRnIVNiUF3eD8ey5bvrrT0z/1Ywi7n5WTcWOkj3TIEvmIjKN/iJH7KCrUO
QdLlz/cZeiKGQWfoVaTQX9ThkB+jZ8xshtnJJwRacQDfgctnY7Owa+S50iR9Z2kAId7+IycnprN6
gGcKjaHlvX3YIAfBKEJlfjXdfU1B49JubCHkjjqEnx1jTNI2OROCAukZ+qjHEJl2yArKdpw4J+zq
zV+t2wVf3f1DesopiHeSQVAlCa/VAL4xNIPZMjrOTw6HDgNWUOPGS7St/6RffaiTiAPhbN2vkhLQ
55dynHhBpcQHEZLN+jq7IEIq6PEHC+MycBbUqFKoN7QAj2r89q2VgDTU250ONhNii4vGkQ4u7w6Z
NjcModcyiTACn7Wx/79ZliLF4QSNc4tlYzLXg7RnL6cXsI1KV8Qoebmbd3sC1KNCoCICCQ6N1rEE
dfrzcNSNU53QM9Ozei14YaMHsPWYdD9qpqOGB/4iiOdqXF1mLA6ZZyJU8cFMev/yQB9IpmFp4NEK
Qm/uaajpCU4A24gNxhOQxHfL9s7qLSr1dDcu+U8OcQeD7SYINnqo9hxDCzJtvMBQuRqrgarF66f9
Jnu2+6M7UUTjuEoNlgjNs+9pUbXTQ74dpYol1IOYC1tSAgfMPs5/mD5eTAFipUAP2gKOkcJij5Py
0zPndEtP4HuwzXvhIQ0Eb6uweWTnUR0cp/aK2T6VTKTxYpAIVeW3TavFr0TASGT8maox1koCpilq
awFgHPl3x5k2jxTNrjsLWyLBc7O7CcUyzdHFeR+wJFkVjqNqEPtt8kguBhnOsM6mR8GlpPtfzh3W
Sb7ENFHhzjdOueOs3H1EaQ5A7nND3tUjHyvM9hE8+Gw/Oh1qa3SUdUTx0rZ7/k+SHJzYPRz0yLsd
nOiPqObwAs0eKNQYi1X8m/EI5eiP+mmGD96nx+2nKmwBa6i5pr/+RdFtNdjLWlqEfZi7NjjQE/i+
7+KbO5kBTWUFiRFCJq+ApriNuicfDAmttqpVsYBw1KNwjvgN/vknOI2htyj64KkkVIbTCOuL4qP8
Kgrm+ISonX8FyrO07LzSoOW1sTtd0DO0c5Qy8NWC/dBNbf9bLIQ0On8khTjK8sLmOkLwikh1QFlJ
lZM7U2cHvxsVQZRAIm9t3Leu9VR4hK+xQ7c4svHADpTx6QQXBkjcZZB7pNo5MS/7RKJ8XT5hFt4K
Kznva3/IdZ07OxLunrwNX/XkD/nTL7RtzhRVGf6fr7c9qX3xxfdOAeAK3yW43ktNsWmrxS5zYThf
tU7iRTtHNdNhOr+W4OWeu5MaueG50wCHMmap0nKF7zcUh9SQKQ87kJfqFiO4j2np5ZZTCc7pd6rk
hQEOzb2tyRmKYYS5PDjwrob+s/6QiYzcOk0fvZ1wbnwC8f9HYQXO1Y/1RDuBxbPaK2PRhaUVdKju
ywr18MO5he+AMUCPADVRiZUVRFgrK589uA0nNZWfkBydp02go7anzgmQcbFQSMcTEzdUelZCfBTd
0n3ut3rMvkK+XT0CPBMXgTzX9my/vS51CjXpZkINESPnR1oQMvZy0MyEMo8VfgBB+4Sh0NfcnzYd
MhphJZM4D4Zm9YYzzA9z1Y4ViU/cIzBvnH9609mkgcdHn1RHV8TuawAe+E6t17rwYlwQlbXKREMI
41Px2jcHL76+FL3aNmCSwqjjf03SwTBkwhV76DetLcAK9cPjgAbftiAhE8IhX3lneSy/NGvhfR23
aSoMyU9NBfcbGmKhUfroyhonRIB3YlLTXuGd3AbDN1fPU3xjhlRzW6A2rwWq0gwnw4LFwHmd68nU
pqAtEp/is0HwTpjSuHxSL2M6N8AN7tCRXJbcbD6T56m9Hbn5JN4oQrjG2WSVHbzYtGTPjPTvh9FK
WcblSWUqmT7US0ufYL/qw9CmeKqf7/aflGYhY00Bm5xse2HkQ3RktWYfnqU6IZuhNYRIRbqk3rMZ
ncMXLcCfBQasrg1EVFTIX6TW+gOM4GX7GABW1onhO4dxZMSwKBD9TtHD2KvSCUajv/ObEQeRkgjz
4vWkrSRF9DCjF6fSmPxTBaC9UoFEsSrS+Se0BbGyvtMMGPLwT0uw8dlK/nP96+8l9vwK9VzBPwxY
XE3bvEdaiaQFRPpqMGESFfibi3bLDsadJ3+2OKRGNtkPq0R8i9tHPwpnZylF7ONT2ByHEBfDRNch
+j/7ipB1CqLPBaLSdOjf96EAgP+qds+CSW0Hhsb5VYwW7m1tT8xjhHiqkOjzIR5oaa66F4YH5865
WJ8L65XfNwhINzo9yvUZ54ekHaEnyXRbWvlhxgyWgqTq7PR3Fu71mRtLxGsbeEfqMcxBol0n6qQT
DrxstXP8b+JyfDvPJNVrD1QRE+cQfP2/KNoqPXga+IrzmRNLJkA3exbuell76Mv9jcDCoEQSw1FT
9dxX8T/3sxFZIKUfSCiQ4zoERnUk1RVbtSX8lzd9SVCpbPpzzl7KKEwSOlFFuHFcikvaXLMsfPwS
LpiP9bDeBsvan1KCxknzCPFccTyC3ai+A0U8T56sWjqguIBAaeeC8SE3dLOPw2FFmMrxe9OdHplz
dk+Dz9pWs2tU53gFy6Jw68DNf+LmtL+/oU5UGdhkIhrwxzWIYwenacllpG2oSRTIYalFHYpFQkt5
tCVPF1Q0K5j9xK4pUstv7HeZgtbBNQVS8sQjaxStv//jCFP5i4HUDjP88Pew2rjygK9p/nqJ/y2X
B+Z7/v9SdMmMU+9oxS2D2AoFo0s6cYCt/YvoZhJgdnVNW/rijioMML2/vz7t2NJkUsKK3GfoF2P3
tTss/smB9J+60NWWCtPHy9niPbRnj03VySjwFKMM9cKIhgh60Iq7O9VgiOImj/i0tTKDcCEeyhV8
ZTcw0/LopzBkvCkrs68nFexpbhk481YS9xJtbl8Khbj6XH/2E2BAu3R91Mx4NduNe95YMpYD6PJb
22kd1XQbfVD1pFW7oheFyUzsBT1vUAFU/roa3JThSFq+8lXfTWxgsJHC6tUR9GZMU+Xl3iO+Mfmr
mZgdg18RFVq8/YgafSyT+uWTVbMkgKwEdec+VtsR3XCc/l8WsCOvdheEd/br8FO40cnF6imc3lEd
W0Axva04ZKQysta3LZGLYhc8WTWus8R57EaFx9bZ0A0Vfuk10+01iF99pLJsOwStvvCLlmorC58J
oR/N1CuzujiPmWumr0HtVvong3NQ1JUfiZe0GrjtpdLZpXhnwzp1YIG0j3lIuhLFlns8yWIKEONm
zeO6CIIH2NH1MpDFn3zFqNStlwadq0O4DaAE7Whdcq7tol5FGLxcRZA95HdPagheX6nieRT1UPob
bxPvnp7Fqsjqfh3JUpwgD6fSId8KT6zPUmKahCqg/bAtIJJyCmkVTiZBoI58k68n/FK1YLQjxjUV
AengornHzN6X1Yrw/2sbW0288kBDzab02r3E5UeitOPv2z5EdjBrjf9S/WvXXOVKUr2iwFRzDEUo
7Jlt18P53zTRXmilSh01nVgNb49MDooLB9Z0UsMCQYhNM2uer3Yo/LzXQ/d4fP7pVc/7MMlJCm+q
7kqvlTRaZESqdmLY8WEwyeBtn24hvX0XzQrQJTfYENGk/zNDvxKosRsBuioUE1y64HZXADNhgv4Y
MIfq7miWOaovmltrLsiKFsmsfmMIZ6545+Ie3IllpY5LBpUDutOcuy6S8pXbPqnHA56hmLdRk5NB
EqJPrcgS+05G1O1KDcWLXFkt8wQlPM6Deg5RC9uPb/OrCnM6G6tbeoHGCrqSoMZRz9ZQ86VfCIOv
sPT3Nzv5Vbbk1WUowTydGnL+Zgge/uvxMZTy7XClgEoC8q8mwyHuSKMYFiFeldcbkI/OhxF8ZoXV
mEhS02ariPhSKJ0qYepFRf5lgj641C063Vh8WyoRUI5Zrpn19m97aPfnrYtK783+Dy0inBm6ZaUv
82dl43Dv8vbnGtA7W6F1cV/L979mqceYScoTZeCsab5kcowpVKhAewsA3Yq9R/XY972WeoflYwZN
Qo16K+d8gOTaM/ynJxiSWui/LeNTiK5V1A0mt4EMIIxqRam/NuQFwx5zPZuweqYrc38ppdeI9kOl
Mn6jEl78/OYQJcDpw9cLMvhoBQgnxZ6/G7DfgWTNUg/rEDYXGqpvWUnIpioebrwK2FxXZspdabHt
JuJ7nk/IlJfmkSNc3dIicS6OvBd/BoPLTKaYPoRwURm5GjYlM6cnpF8xFDdf6Oh2WR8If5papwI6
1dW90JCJqEieQgYoQMBOJUHpwhW9ai7EAjba2ezK+EVtRdUPZu/4XytFb6zYTqIUOkk/1/rhrdgh
J7H5gcuH6YZg7TU0Ms8HQh2NZCYBlTIGOENaeyDapdSEVLH8RvEo6HC7mTU1hORjlcqo9KtPXm2F
HS8ePxsCi3kccIVUgtvU3LxP4Q5nYa7vTkrEzfBfU+uTr0hTwYd+e6Q00JJZbrQcitT8+T2crZtr
E8ITdnqtkHRSDLA54vO34QtHwS01mZNZyyqMbSm+mHTFsBzbSuZZD+WC/RTLJPSoiI+Ed9aXPoBM
Ov5JT4iyKHDD2yAOYq68qCEfA1sgJ7tKPvJNABAWHIqijFuKRLkxmfTUKaQrfZHmq9nZf/3waUT4
fbayOHQ0g2QJ5Czo3s/72idM7YTmxGh5Q7iOF6J30XDNAexLVMHpmi28GmqWiM3f5FSjbQNWb0k7
OM8h4fIPCtd4wvGG70LY3eSMxQRPaUaPj+HIVZHhH/1aBE2XCy+OdtXwtEAqfLXVHZAssgn/sPd1
Fwi8+QSBan21cFQgIj9H201+NrpRfGpWgyK21pgWq3ATRSci3gugthtLI7Oe+sYXBqq5sOreN9yI
6aGFOw8ODFiVNh1+inkHzYiO3H/lCgnRxacwo3qhsTxbUcyF3AaK+ch9mJHWS6QVepT3cr7JiqFp
v/xwfXWJ8KyKklXJNc96jUNPM90Vj2JLoJQ7I72uS85K8CbyX6Nip0RbEmCK/ZN+JxggdCo/Egc+
SRP3G3W2N6taciA7Ghqxs13RLSZfPqNs+d+y6bJdpkEzAK4ANz0Nwg6Lqibf9r6tdxuWHP2CwmQ2
VnifYSQ7TAM6usskzlGOf+ieHeErkMrRJjtXxZP93IE/7Tzur/JFHj3WIN60lug4LWSiNX4vtBgJ
VmQkJvsavomi5Dv2eWahDPGwBeXSxd8usXbeNs8D9a3drNhNZ6LOxwOq3VAu59gb2pzGXq5GAt75
/qukj9EpMfs8b0oqSMPoIk5O0XE3q/YACu/BlAfkAd0sQNW7DElpN8Tr+wqyxJ6vXHS5p6UnzIcP
Kkfsk3nY8d40dJt/z78O2tECw5CyzzEOqC2sMLjkkgB+oDUUMxZHSxMf9y6d+OSOVqGBBCOlk4My
z2YHHtlCdKp00BpEVEu0RqYUacthQCqUlDY7LsJHaU3wvORIgDoAlw+a9DqEGCqPU3MYnv0xRSCg
X5OQ+ZY4BzHv60+G2N9HKxrpptLedrjQPgAA9PSmEHY3dp5Y+PE6xHdTHCTLnIcN/wXmxYpxEMhw
mlsE8ITvQPgtuawvUxP1Lk7zI4jhEU/B0y55dA4jwIuaJpJe2J3g7ojL3iQag6had4Ij/P6+ahX7
ggN3S/+1nC7y71jt4tyk3PMk4HbpuqXcoLNk7WbWOSMA7ECchcnhtHRF8qlEe9IHiWavK7vPbtq7
yajZyGvlQ+N+EJTfv+ROsX+JX0Axtr0Gsapc8wgeMFLO31B81yPT1kBfR/5w6HoSFmxEEsJuwPiT
pH9YO32FfOYz0/0shD85R5eApSdo0hjO7Czjt6FFF3qezUsS+NAlWiu+L+7X2U61XGSsgZto2HRb
Qgv2UO4A1qCfIP2+9Xj04hEihJGdutPF19iNnROhR9iSGGDIiRV4JuDKrlQEvb5F1T696GgIuml9
2BO22oIDyk7Pr3mh1OT0HBw+2fzNCzRZ0UdeYUAL9MZ8Nj+C8iYa44MB31SCIpaYfJKx4mvhOAYo
hRdFNada8KNo8zsQGeobJi2VBOSSWbTS70RBYGHzYx80NbYJQV/QtOpFQNNqVtk9giqI5jEgXF2m
lw9xf/++xUDDcKY6kCDhkq0tgyl9Awx8K5L0iy0rnGwfghGUwT89qPdY4Hv9c2JCZ25yDMccbiv8
WrE1gS61fMJSm8WBEDMHHCgBbviCNVvPPJ3qSRk6Cq7nv0mGTh0wrVfxplsOsb7esLbzH3Lg9136
Dml1/99HrBZvkTjqQ/Vugd5a0SeQVVwQMXn0lUQH3G27jaC94lsKzLW39EWbmYymadk7Khxqndoe
z4ECyCb2Vv0xPrS2RX8og7HuTyoLVIb7zzi4g3AIxIvKrZlCUNsBl4I5PPb+QhxV8S/rnqu18P6t
uGrABuB2c/euxzAyIvMQtPBLGkjiAqL4LIIToWyiCwCeZD8ezi2ac8xZ8s7is6A6C0DvlIZGGTA9
Nm1/IPeyKO4Ffvy4ncVtFLYVzTo/5U9G8/i5EnHroPSVOd1U+R8qUfSgpObrF9d0tNcgTVwjwIOp
CrHwrSzN2OozbW9raXpw+Eb9qztQQDfpZW+x0td3/tJqlAcr3ShsZZjHSK+j3DuO/kNHnlE0yopi
NfwjdAqIkIVWHIqiDqJ6Uc+PGobrfN/O2h5aI1m5qAAiy2U+fQO0gQUm8z+p+yuBrIMJlrbXWyCB
AddGDqN8yKF5+OQHs/bU9C0SxpgexSaFSAcEb27s1eJb77gQ73FfjTj4k6HkBKk6vzeYKmz2Dclx
yoZAGi+PvJ3LY/VAbh5HLDOQWgCfbPT6QXZtedcwq9l38ezzOwbWSuD+51p6SmcGgxMI4KZ7VmK7
TDVd3PUhnIZkYwd2DDaay+swNPYXYUj5y6TqS7UuZOaQArY6WgZtgSCKQF0FTyqPxh8VRbyOP8IA
7Isi8voBi3cO/eC40w9bYC48FnT3tYd2mggxbFGQjN27LEz6QbSbtDRWufL1/lV8wb6Ia2lH7yLN
wYqz6d/M+6a/Zosd78rWLynmvH5mFvYsZBS6LJLHEfpeH8sVecPpNbwn2nG5e8ZKqzKQg9Nvpn4t
xuOBQe45ekcEJfGxvwWCmojGq28AqY+WO+vhG4Uu/KVYLTCktwyjqA6Dq2+1qp/SdVR3ZXsX3O4g
VWs8cUwWVjLGwxDBkgZAmTsnNHj7+kEqai9iZMLfsW4HWdZTMEvIqEwgEUPmPGkqKo6SCUdLSFxj
iR1ow6/nB9tRFJ/IGopUl10bin+tlU6MYluU3CQSITflv3aKqNo66Gwt+Oi1tkT55PMiQu6NrdzJ
x0KDDOIYkg/UfR5DsxbOOoFwnubeaNQsHuOafcy/K8BrRnNamwIUCB14i1iDrp7nCkD7GLH3rpKw
Gd3oTYQJDtg2iE6LVu6zRLPYNqu1+Eg7tnHPM2boBgX3JX6zcYCAuhnQxkoRe+DLYz+4tea36MCc
sJNFgVjLccEKb6BE0mJ4pqVvST3v29/pM5w1nEyXFWVBwY8SvaFW5HvUzGcNWblbIfnxefEpw54H
ZQvSd9KcabmV3r7zMPqtRZp3Gi5HYLyb/guOKZcEgZUhOIVdhGnAmTuy8U23BSAbeUfXnxh73+iH
tB9NUKylGsv2/WKSk0Z/Zzkf36HZ4D+guQV+PYCsg61iyoDJLLpAx+XEbrpc+LGpUfxpZYryp9d9
W/+xS1Wq1Q8b7H0GCps25paXV7L5yeT4z7GrC43lVvUZTwL5kvia4OKWFAupjDUwdKrcRy6M+GR2
/Yd4TB1aFDXPDeHgCJcAf+oZxAc1PKu2iRZSWTYRcpSK+rmDuZg7xvp16fL0nfhNerDiHd6GLCC9
93e1ivq6Z6SjQAb0b+ceXxLb++1DttmB7WCAT7f4etLbJ36+A2297gJ3p0KDD7Unq9QN1DwfoylM
7I/l4cYoGKthO6Vc5Deq6F6ktgYK+XqvGJOKkC0/FY7n5NtoNhZyMB/nrCQH9tDat1AYky7VjqgQ
Drm8g0zxR3mTxq8aOJWuaYlEGSj08M9ccPfTI4488mSCkArht36jMRs9lgl7StuddcRLG4cilFUl
fpM5Qa4FBj0JSP5rwILCq4rlrQxxCTatISWgd6Ct5JcRCmF3Tc7Fup6GC0juplQMoBtN1KmIgqIN
U+0oCCyT5sj/4aYhK+/UaQzXRpkmY5zM9HNNv5D8oluR2yDIfuJUiX6LhMZ8KtMV+QIM67BZPV/s
TV0VgDeBtdXO+MHN96qgM07tOfT5OJh35NNWQ+Z4cyfqMIy7M5+KQRn/apXEUPWtJ3ashQQQ38Xb
fbwlonv3fUWqy1SjfM/1+in4ggTIE+x8h0KohKIEgaLOtKhpvttkNmKTJl/xeypklXUj4WlkZ5Y2
MzdjDJ2nfTjwz+9C68HKzNcKOCikEIAxvqOpkZx2AtIJh0hAPwvdPqorWCiTmCmW1TCFRd9bYTE2
9C0UwaG+suXT+/2xWj+vpL/F/4yO0hw8Mf16KuxMDVNfuE7aSZg3R2i3rDGfbDYUExbss4ZCkMbd
FIUpRoRRGnuGqUJzxYnCJ8E6jBVXCSV1NYN7uhuz2ta4FmwqvkqB/2O3d7guVQTRH1diu/hm9cFV
hr/bTKW7t28jeXHOf7MSMit5BtO9ac5tRkrzJORp7EG2VPXA95J2N1xo6Q1hNqd4lS9Ehaqi24BV
TAiUjiGT6ulrj5ySm/b5tmA8+rVg+VM0cEk2rReU0FCbMRiWG2MwY/iwSst55Cu7DcAvEMjnoR+g
YFiIOZi/VWZxbF6XPU1uWx9HZC5JMqd+40fs/ig7i1MtFNLm08Q6n1wiiLOi5EOBceqevng8NgZM
ROoFR3zhxKFEWHd/qiV/0FpEFsM/0qm2ZieENzVzzwVTQvM4WuedoTJqByMojITvELL1W4b8V2pQ
IfkSpBPmsCAsyh6bVEQL0mCOVh5+koyBHVEir61UZM/5s+3aNDowCJbvBkZHJTRupB4Vx11cfb9h
4v9z0gNLyEUTzPjBPCco7w0UmXZSiito8TQOn98JmW4RlawLryzWQzk6xvp40lQ/OgpAFbeOY1ir
yxByi9SHDMV1i1JZ0MwNE3RbR4aoqrqm1pefAEOceJcle6C0BVVs1txVJFETStnC6HZmAPNU6wPB
wnL6WMXqqQOsToWRnvhh1S1e5+Mju3f8gE7JQEjQYH6JNpU3lzS6Lvlx1caFGklgQV3MgvTr2roU
Dj1O7fZOwFOwyIrvZM/MxsovrLxi5Sv8ywalfa6dZnh9WZj8kjHnJ9w0NO93U8QWowiYSbzUAHHe
ee5f59/AmjZ6APgLOIat92eMg6fotgR0rVUHksoMdg3JHIDDedXUcc+YqeEvPz07l5obH6MVEu30
em/J2wCdEgYfd5c12RgxOA3XPd3VwWSyye9Z68OMtu7yDHiiPwPsPx9Kmm62WjUuGHrQmCFPemr3
wHH5VJ+XIVRLY691/OtPU3Gv40N0EaOUqGNpx8RYe0TFWCyhxaZYGCC2dMYR771UVulRO7Cu2NKJ
n0U4CSzHnqi9x+67fKFihcqfkm5xWiv9X0J7eDat5Q7PwLLsZoe0VaS/yMI4Cu9/Vn2U4IM1KOjk
rKAtjfeTnnkB+788eFuSyuzAyhOdXAk2eFESw1d+qJPtR/Od3aM+y8JzppM12mtI8zSR03+z0KJY
ycGDauHf1FBXDVCb+dCVCQa1SR8a5szLsWx30OX6GeRPnwY0M6T0xrnYP0pObE6TnlrtR2MwlRNQ
vgUcBpq9KsyRDxqu381uc3i6L9pJevvzUwDbEMP6HNT0XH7A8EZdaZjPMkMYkGExL5Flh1bJxzOH
+XHFqTGWB0+HgOIM5cQ05pUrp/KzIS1m8nji0o6TlNe6OjbwM1g+1d2XOgbbayz060ykqe8GxHqz
Cnazz0d+wVo5nFpvJD6pUaXqpfzeytgT+nOoh+L2SropNaNtCvb06uwzCWsN9x7QlB9rc58b9h+m
v8Thg6GISqaCNrRF6z+Ht+zUI1TJjh+yc9dgCNNXWCqDv/qFEtbDRw7uHT5iIpBLItyiVjWB9TJl
dHFddPTcwariy3mn314dF7vscy29yX4oz9sZ4r/rm2aKzIT+0olnMtyb6PzXUkeEa9Yapi78nEWX
rHt7PUokue+kTkLAh4aPVTdQ1peWz68FinsFvZQi40KC48ITelrBYV/G8dqpcNResNDC84bxltMh
pTACWEWGrFvmRsJTB8JTPCVgCk3mVQ2i3QxIgeFVIgM8UQxd1n2mWLXDpPmIz47GyKGkwQIqr+pR
PNw5VqYRiE53kwfe1JYWzj+Dw9Ya1ffJdhUFhEV9lTbY7q+xhjyZxtHYKAI2Wwp7O2jVwqOxfDMU
YSPVTRJipoJMEiJ4XDkjJZtuTwD/aN3tyDcbu4fKsjbh62dutyxXHj2HpbN6kcnRWCeca6H69bPH
wVTGb/nHY7GNBI81QGIuISfzaMqFocOm2yoTuzvUQ8ihqNx5i/v2KRfqCUNXUAOyUGWNvgH5CcNi
6yRN96XZFxP6fHyfQSJOsLaCcN4/I0ATL3QS+F+YScEP2z6bnoj7DHNMkkdTf8ixfbJMCOdHvaOr
n17WcaozYaNP7i1/84IVhkLN1JlqvAAsXhmWpmQN43EZwC1y85b1afu2Pd6SKVNzMHuWjeEKG9l7
e7YHP0F4D9XEgDTl4SK7HsRgVpxAc5ocW3MUfPBiux1mODr4chS1QVj6GXAYGt09I4eIQe/BZ0/Z
+TEolyszX+Rrhyrx9n941q8Uon8Q5u/Q9P7ySY594Kvphd3AwQAkZxzrUsm8ht0AidZ2Wt5b8TpR
u9mok/cW0rjd0FcZlVpe6R17kkes2B25EKPt+08K7gd0owpq74N9ZxQr/LkkhXqF5M/BZ7kZauUP
dFNeNGKDl+jKIykTd4pd69F5zicmVbfGE0dMnmQ2v9k820SKY6au/9FvqE+NRq+hSzV55j1THNYc
anJAIJD+xqk6rBdIDuXlF83A501A5x58f41RrM/lpwBWeESX8E32CAcK/An7dCGtg3f+jh53blny
vANkDQDgXgwdQtxKBTCR10+7JMCWHeyJukew9Njpv61vA/tzbqmSQyqlfDG00Yy2KTrpc2zgJE5E
3cyNAfjvYsqdPwmSSrwCCulhKk6AdPt078+u+e+PlvSdetEC/DvWYBrB8dxYpbo9tZVnbVPe5LUX
l5EcK8tCtJtx/QeK6EwOgu6o6q8S83PGfdLFhOX29czfQU4F8y18rEfXtmWoUmAtmwwPH2rZq04L
ujk0nBa2isG1dD54qPnUShfCTFj/GN7piU5TpebGxze1xSmNs3CRoK9fLAQU5u9dmgi6tlAsMqtT
XZuDmGKptjrXMK2ECH6myzUS6GMyIdh0avUX3mtzZjM/WJ/6lEewlqfqJkGWAvlBGlKa+DboQNNn
DO731RzQcAK5BVIIw7r1ZufDgYz8j/MjSHLQFnHkJtr63rGFmrHbgkD90mdVaNgZI6o7Rb9MFbI5
iHeMHWyIXiBrOuvvnxt1yWthcTajNwCcm8LI5UgNUNeTb+VH7crvQ1VcJPCo2PIo++4DWxU9Rgrv
1Spn2gsdjXICv9ArsxXHXfIYAxlWv4i/zIOX3VMfabDEA4XOHXPr+YJc22CgaS70TF5ls18r2WrG
UUujdzPFFmVK4zrNDoM7sdJXxRvuvYgL28Nt1Gis22+2dTbqgjHaJ8FANQCPzK+DytcPZKJ2C0uF
zG8coXSlX1G4d+ttYNLLhDjYP9e+bnEbC/qFM0PHIWl+Qf2XRNBK4WjiXT7B4j/UIuxIZm9KcDgG
OXrXRfB4XrJUiJpj39SoZlCCoN/SkZcNVO7gyJAYi18u0z+A723+yO3r8c/EwwLz97Y/4urOiOAR
9Bw8fHTbZsB6SbBUS9nKEnIAeCgmIlkuTZZI2+wJt8U+AxXhjGij2uGIaAm8cmNSN2VLaqbf0a8g
8ndB/yQ4f5YRVSJjylrjPv57Y34vRZ/XRANc6JGmrIDLrtbwCH3zfDk5kXMwDfpI9j6vvWCDM3Nn
sf1vwQGp49maavjjg700OTK/8Ngw2ytMFyC3hMDDLlwsF2zVUqtHkbhPOHp1At9YPsbbxdC9CbSK
HhjiNslbmcrS/Uf+tGZ6cEw2gFU7lIocYmvlUQGQl8DRw+/6Ifvgsu16e1vUbp6oS7h2JF2LCs5D
DwTYPL+9SOTT+Wo9jBheRVTatzHgtS6MX9b8vmOPsU+Wj23r9xsygdj+r9yeNWbXSSCmCY2p1plR
vOet1zwysJm0807Pi4yNMSnEHcam9xq8UdtWFNsJ2nW9PMzf1sHNCoaUjMeaq1m8k6lVDCIzHDp9
cfGAq/Z4NDmW7ULhQbsDR721lQ7kJ6oh0q3TRoQ+LZvZBhCCXHUmD92pTY9KhJZLxtpG1LqedJyE
kBwXFp8C2FcdSCDXKVP3vdkaUZaqbYZ4LMeG0RaaGrIxAV2/5c0JLgzVxSCk7oJ3nUX4mP+dWF8x
s1geux2L/iGeQVrVI9zEKJQdS5wH5JHnCnAn/jZFYf+HFNYsPFl3t3kcfgpiO1+aMmiO4Cv+Q/V8
b83Am0vB5oTG+OHFo2YZFLTytozgfqZ63WJ+UrhIxegbKPb+hOKLjd4S7Bq2NhQNlQ42+uVupzzB
1vKkZLHxLF1rkBrPAgxx9vvGZwUdlCzEsFba0nPoxYDxbnA260dSCnJ723GWCioVXadMVBzgAzpf
GSSm7CS5U0sNo953VwJotgmxF3WxPoAm3BGksl6cTZ6iYGdM+ZYZwOi2Trkjgm2Raw1kNRb/XK4h
OTPDki8uFuD/NLnieX7F/LzH8OH057R4xW0uQXQ67uFFpNZof5i9SOB3KllICnqRLURb+ovKASrd
hni023HFuDd/48PJ0MxIvt5ESFtld+cNTArnxqMUH0nbM/O2gGnMFCa0/uEgp4jH1NNKCNoroGKN
sf7LlKPG79Z81kIXlkNs6dUukbxSNRmIWq08LqR9j4XHEWz3eS4LudSIGQZf4jsb3mGKE71CC+7R
u3Bv352+DGkWsaClScMUkqxq4tpdWD39U1BxJRqNjDIVqjHSatMQ0zMo5JTZrh3Vang8OZqPFAVb
5dnV2cybU19Ulr/KTz+zXY/bQEo7upA+m8oxZdfna/+XIvuIL3UavXUXthpFJJTU2i6ZPjkSW3mc
9qWLfg70x9wVQjNq08beYospq2ggAumf44QtqYvkr3SnRQPZjlqGzB94yKDPZDyqqcGgfOATVSPM
uQcmlGTyVKigxvW9OE7bTcKy5oCTjWKef4aSLaecHIkES9Dly0I92WTVZakXILFh74zAm/U7ZMWs
CvUh6qyZ3KsIs5m1o/H7/sCUqEnr107uc1t4SZ64zWS/RIcFkIEsJcLJazh53vRCuCmNtAd39uE6
H9XPcbtqnsouVd0ZhDHCLzd+nieatg1v5D0tf3M9bMxYXIRGzr5WIOWt5UdLaY9xMxAbomCl3Bfu
ed9EBOdKNFAZ3XdOoYXNmOCaZpbmDNf/mbjxEq1DqCNS5zphxnlN7dPJpodtiEktd3HMvSjYPcg5
w6uPpoedwhZs6HwTn6iETp0SQ9HS9QD+MPgcvyMsvfD6jTQ4j49mVSu5TsMqAj3+YIiQwbIYze/t
knm9NtXC7ZFWdbjpaoloW9BX/YJKtt+ddkdJBjyxuj07nAtfV9yBGAPBeF7biIgBi593/CWqh7bm
YIz+6fofSrtAGoGDY/DUnq9QXdHhz11S2EJffVmClexT5jtNNUYnJdzfSsd2E8IT21wCHQCQP2Mu
nXK4gCyWe5+6Kx/RboV/d59Lh4kwJrkbrsdiobk/I2OuAx3L2KtSYT56fx0TMeACuBcl6958V0Rw
BxG+84IoAjPhkCBQ/F3eG/g/2I4cTCd5QQdkJ2RSKhmBN6tv4i13Uw7EweSasCTm0juRPN1AeuSY
3fUbRbAFHTXEbfnzskY+zxWC3IWywW2GVxvN1Rw08KGAEqYZALTJkBK/8T3nf4GfwPiWcKK5/UrL
S/eGUCARRQZcuYL2Z2tnJd91mbDl8oWRRQE9DF1XT3kZDH/fjfalh8CsHh2T//HMXAoaBE8jaU56
LVRKjZJxyt4eWMQniLghEQhzlE9lzMC1TCvjoxBOduC1uvS0nrS8IQG4zllTACwJ9AviU4KXMj4X
HCZRErE82fCEaoLGo7Vy6EjkiqBD7Hxg3XcO4jaFZpcdXeJer4rxwunRa38f2uQT5TjiuW1wjizC
K++/Y8Lb2SoXrEuUkkvD6UoVwHawKdlvLTQZBpFfPl3c6aWzRiEarJudQuQZtklOO5TtdBDUavq8
aMutTcqoqCVwbqMSLaQY8my0jKTaUxp4pa3Rg/SnwYs4MDscKFVBwn4LNDNKKwzRL/+OjFNB5lfF
lP6vbjA0R0W3nAFy6oce+y+66CkBCZBjgo6PJrYW/eo5fTvdeKHzurR3DlF3c1hMvMxEWEnNQ13/
sCAJ+Xs+jW32vB/j37BlFRi25DKCgw4e+NtR0UJv9HBqMLheYYKJu3dEfn8EkAfM7HVYitGpDpQf
FqD1fDSAmdIv+FqmRjBS46vfuUJoBpB6fRcQpPOjFrqXRKgegxxjlCkcR/OqI1w5V7fBgaHdFu0v
tU1zGH09y5O3XWqj0yuPhRklM/3WXk1vfKfLeLWntEspRUuzj0jhH9G8mpMLuaquwO6GsR5sh578
pXS6oU5OWQ6/4/GB/yvQBQV7caUjwPhsVj3J2MiqnroajPW+ljBGipVeyHbBQC6jVS2CaaPVv34L
myoD6N29VghaQ3ItrG9aLq0WL48cnu9Jro1UwhwTaPhrtTlbU012j9c86SnvBkzJKLaPWuoO/OYn
c53YmGMhATvQLMpexXx2n6FLHojKfe1By1XVY350yU5oIurB7UKxUKoKC/j3pYA5zZLL1uNSRUtP
tmCvxKYDGiOa7sjdbwWqR2XdwIPrw708FS/akXhap7dAo9iQOi2ilCmWr5uWN7CJIQoSIM4hNniO
FZhkZTPEmTe2bIUoegJDeYEAvPeJLOtZ2nghL0KbUh/0pkVjzdN9NuFvbSoTYSQtdBiC4J7T+m/D
MwbI+/jBXIxSAG/f/mnScoDq+Mzgm6VZmwRjVyFxDf2ZYt55kBSMBbQSO+Oo/Z4fKUuOMJbI3kkP
mul8dJ8sMX8NK6GLxSXTCRuYg7qeuTgNFfIxJhYP+jtPoa5x0nknz8jR2RtBnkzxGdhzrwD2ABSK
NBEIhQVvZ2K+yxDGu7+OQyfuWn88JvI2jZXfPRa+70vJZbZNpwjFMYmzsIqcBqPbjpyOB/pm7bAT
HuL3q57/KJb7Aam7zLmhw4+iQYBPJyifdhm1+lBpUoVzH88LjY1tYlZanCkjgyykg1FyOVorftap
e3VENf333kqg9pgChkCRhnLIAjFp+LXELaLq9NKbq/rz0QkywCPENHmVy22oC5c2X4+CyrbC5Zr5
vfBWgjp2EBYTBH86LT6s9MzYO2ThpxvgHuPGUsSFvi36rIgTmvpmMBpnHXaYQSrp4PYG1fV6OhII
HISFd6W5GvqtpDyOoeQ3NM7NGj81h3A8SJcM7SJJhCqKgYS6JI3nAGafFjUOdVBHF0efm9Mi9ew8
Ot5OPvQNVBKGhkAHTkM5owBsPf8R+h1DeJ3gDaYGOrmtmpbLsjRUm7DEYB9ph6mQlKeb6KtFcclB
FGwgIw0ipd1VbsU7sllWAdzXNLbexU3CunD3TW2itWq/b3kbvYtPW5Lt08VzrJ2bLDsinUjNmS+W
Ag2FWsgyid1CgefV6rWRfWDS0szLQtI4JaDi7ESBzFf/08MUvhciLE5vFELLLQ9Tzaa1EchV4wQy
swxkt5wLSRtx5+VaZmIDd73AnGKqfznDAzNQsPECdP+5ukYdTuH77en50lYColHNTxVujSrYmL3e
Y2JEe2kOQ+1u/zzntHHXNvEt7WBI99Evx7SyAkSAOIQtzvQuxqOc67VnCb0039ufKglsd3UVxWWf
4AArZyQQP53a2WfXVM3A1pa3aOQmyU9P+STMlF1HNiEB4zgthmDYs9Skq/wZ7X4uizmU0LQn40F+
7jrGoVM2dFWPj6YzjS+A1ArWYEe+XLBp0kVvJnONqluRQ+11vNoPiVKcrbhdLhGMgkshhzpWmM7g
tclPFJYfwPNrrYwEiNW71c87EHAYLjCqBIxHSh/bxrEhqPfMibSxa8AFnIFmp58hKVCBFnhO5Zq4
QZGmiINbuvBMdV4HuRaMCrw524OZ+58Cl7BJ6gEBZzdanAJJ/wAg91YyudRIL9e4FUDQGi9H74+E
ebXkGlrFK/BMHwBdJfqZ4afNe64KaB1T4vDWb7WAkjW4RRnsSPvcHUfHicaKfEbhxxouxyHcSdRr
teDBatcMjhioflb5LhF/nQcx8CLI8PwiXdJ5U6yCbyEnKHIZi4CuLu+he7nn1mdSbzR/rm2jX+e+
KqCfXIuAsbBfPk1HZyO440xL9d/S06wo7Sv55nicDpmCZp4Vy0JAOHzons4txYAxCbLW+PpNjTPe
n4VzkOONsLBAZWsxqiHU8i361uuDrchYwwYxtJ8coagbz23bi/ay8ITrfxNVbWPd4L4IH5etfJY2
Ko7GyJ8C7xCOIDbB517lrcQn/uek+x7FXLoqbYnFa/KNf6NumN3ygIROhCCwb8ESFqjBTuQ4FBrr
E7w9pGRupybUjF/bgDa8/3arbxo6bM7zvClddoEaE51E/WVe2NDWUYfzs4GdQ0LX2AP0wui6/KqH
vC66cDSD1MA1Ex5ev4QbNNsTsWIkjQmkoNBNI3HjsfsOtETB8JgWvGW2Jzz7HFc2UCeKbH8oQ9HG
iTyfBga/2zdRR775s3meJ8Dy18M4HOEZmme/0HcjgddH6GGcV2mETcABBTTpgKNzmwxTMHITcU+O
2ftEBs7c/7ZLvYlHAMEs7/+A1y1e4XI/Trsa05Hfq3J3+tP/U0a3NWqpzXgzEdX5AOE4Jl3CeRgl
mHReGA9gD8Q3uUby8n/a9fsTlvJhpPfYvleYJkhi5y1STeYkas+yg3GF1dXFUPjpFd+zKKjg5lf0
y41OwCfz1qaJsJMW32InA4dddi4l3cySgVlG9L2BPRJEhz5tczkMIcYDdbVVZpJJXHXXoQXqdUqf
56gIH20wWEEa+vLHzbrAvhWKio2Tuiwb17qHbFE31RYWEOAnz+X4TrqbsC+Oszm4AQH8ZAggTU6e
dC4iG9VI7WLcLAVEmX0h9x6WZjZZRCh3Nm36xywaYl28cbrzAof3LwyT1/Q8gnH3uxKHWM4M0YFG
MfeCmVzsE1jsA7xEc2rRQ6sPJS7gq376Mez3/6NnjBsunbixEEouUR81f53ZrC//feiVFq7IKXb+
guVarPyuU09ZlveNVK/byEq/uKG3fYm5g40Au3lTajau2tDoxvwFhPzl9kNzzoq2cNP/RWskSRy5
BG2Spse9UE8tBtdd8H7VTaeHxSN9ugLPNJd8jvAIN6gAcqGVMcnLGtJe0JNATd+Z4J1d1+pt6mNn
fic+6q13XlY6LGgwSOl7xsoC+ZpQqLuO5NQUf4wLnVhLj5L84+roSa1hmYKTUANEVxWzO1PnWLWa
9iXPll36a9Pm43sl1Vde7OH0YQSE9qDRbj7Rmbhw04v3aQabhy7IyzncmGue9tUgVC+FHkHlkz71
Oe3Q9josfCXkPTplncZhZ1ROY+RqkI+TTLiCCm2Jy2s0XvefhAMKLHYoIaoZApJQ8kEufc/wWL/v
KanzYZT7vgKDMrIOkKMNcZiozhd0QHOItRHn1fYKtLqBG5lrj/RNaY/IF3i+LqvKKJWuawLxIMmB
YGPHq5wI3GYqqFpkCQH5cs/Y2I/JFsP+UfTlDn9MJ8LlX39HVrhds7JKudUZf62HdeclwuEoexFP
vRWQQxq6zs5COqNDQQXxmDkPE/9uaukJGEoUt/eWivkgq0X2/+3vFC4oYeHmVKkFFDfeOoR2sqNN
a4QwJs2T0/pjmp2Ea3A/GxCTPy6zaQ+RdtAcjZmRdmNPO/NCxIeA6NHdsh+3RPIpwP9okJ8dU0Do
AT3Eez08PMa9l7rrfv+tviVjxWgbA2Vu9gAGxMx7DH5qfQ78PC65IMQ6AVgw+vOfheM3I32MLhAf
m+9OEBUpYNxRLOEw+KDoobMpgal3loLXL8zjuCPIbR7biOrKCV9lMG4s2aUWV64ZgjmBJYVoy0sD
fcwmZHjkpj9kGiW3H2jjqnkZalWrrf2z9ZrtELSkvBzOazHcwgtOI7NYFQj4QW979e/JQkgpQNhK
gDTevBGZSW544p6D5kQ6YAn2qusqjB1nsWV/9Sx9JnZnsl4kuDMUo/n86vfrvCwrKb08QVFJzxls
wm3S1clgKETXZ0V9ZYGVkd1xtAO6eB34l5KEizQ3gRmc/qYRyUI56RDjx8IiNpqtg4AINvC9CHPU
NOb4gDo0hRXQ21nlwQXZlKN+vPeqF1q/atLfmeFS8QA+QqBN5+yOlm4H7aL4KwBGte1OX9pAzXbJ
srW+JboUXff4bRXoQlMKePo7JTZfHfBCXy40el1aMU2rnO9L4ckqOQ08kjV8k/0JWUi3op77xJSl
/Bnp9qwE51KbPke7v9zqkUpG1uzUbariIpClTtsaABVWWa6v7EAyOCeUhRV+KZpkDkIE2K3MJCQT
sbMARSI3RvCovkhJq62jtVrTY/McOZNoz7Ry0XHHjgs+WZXKO+HlxLoDW+f2hFbY4hNGG+mT7aBq
ABqAX7nJMb/JqlCg48VC//qnTRz47ff8B0oiIj/Ze69OycyJmGeZ3VXgnv3Nd+1TKPi8gEReb+In
uI6ciTYBGJl1O56rgz4jaMktfcI5OyFBtN5yIIo6FSh3SZsS6R+HQDToPJAhefq3rHAT2E2TeiiP
SN4HgNqpQErfumk6ztLSmpm6w0J5UqAIbjcc90bSIcpl9Jrz4AzO8zHv8nqlN8cMgaIVlq8jSvnS
Ce/ED/YtP+KyemgP1SwC3P12iPmLKTQZILH2McKxyOHA1ihjfA4kSmSArjt0Et71VBWKPskWQ+W6
zMBnTOms5iJvs08eFGhv7EIH9FSkX+DU6YIIEhkW5mn3f0PoAQhtEjExb1mvZ5bLz+5OM+XdDDhe
lAN+nybHKp2aWTG2ri8hs88zMoKU9/572NN5tJsoKkjqXxHHl1S5bFZ0ZWR852rTk4wLrQq7NYWH
TKWiHxP4Cgsh8xPPOMAAuQ/72vYv1Ew9TRc1FPmgSZ7f5MGztyJLfDDR/lGbKJHJ+s/LCdDR7t0w
MCLN/3ezolGfMiAANQ7QclZ/eI080NlL8oTHia4fWpli1LNTtK75P3TQV2PiRYAC589GOrY0xMzy
qhrjy/7e+GDENKqJyo++q9t69LqvEM55kukVczsivJoJxYHjLw/oBw8HiNYQerwZqXdcf/Aj49XP
vds7e0yyC6JOCXmV/BEtjn1ueMk2rmMMusdqzhdI97U6sBxC7RSF8eSFQW3dBC6FBsx6UNc7PHqZ
gGuFOeHIDyQfwcMcq7qJ8afRfyNktMcMKvWVVdcKko/T/CrvE/+Etm6xEQz3l5jOYQn1HIP+r7+8
m/LKI/egu18DK3jibnNbss8vKaLXyqfKb7nhelhL1fF0zsFs4kjqqadj2oN6VAeKnTZrd71rGFlR
iOgV6K57YfP5BKFaetY4YvsThMxgkw3RQELMjo4D+/oon2hvnYqLlxOCpalthPOsmplIqGBc1BOt
pKLNGFSb2kWGyOmo47jIrTSmAYQh2zWRtFhbLf7gNiB20T06Yn7JAgy4Xpkz4a6Lpua8jsArlREJ
+15Ns4aI1OBVMFbehpv3XxmYAmPzGtV/1eSqa/m8wtLxqHDyH4jumKw0/lYGCshc9iDY2/IcI19W
sW2OYB7Up7scptzvym4vE/fD68EzXLjOvY7dPZwUh+g9NGZzNnj5RZibDSWzS+4zNLfwlk9v1V7y
k29CdOjAKgoy6bZ9YsfzN8bgCqw7YXhJtxtLwU7YHpffAnMz8HCPHEjLj6rf6hwxMiXB8SvDorkh
UpSg4PcE+ns0cidRvTxOo7TGTQZp4PGPoT3puPb8yYxy7gUf3zDA0Or3WJVrSxi3JHcScjtaqPl3
Zfs4v8TpW7nGnQDZ5ssK2vYZ8/OmcHZCSfEmzr7lUJtwIIPtjziYLBdz0eIZnd8HNb/gDIoRoxtk
VrhmC59BJYwHvTtIBYsJYOY3RFQXk7oAKFyA5wmN7cFm9RfaGhb0u3Cn9K1uFk/KwvFh6VbcBli4
/UYTzPX5smZxGOiVVT4uuxOTHl2r5dOVwea+kP3U4IMc9AOiqeEkl00hlCfUKYbEWUrCClxD/b8l
s/4GmgDXDfi/Nw99d+Wq7JJ0NYMzTdxA4Yo6kzbgLkZ26giS+UWoYNz3To8j2ITbKYd1tJVW7HXX
AwtysBhyHVuNO59hoH7H1II9N2Mv1WynGRmYkcY+OpRt09Gpbb8bIfEyIyY67xfgdMgfiw61/FF0
XidFHexDOSyDcg6gNdYF2Aqu5SNXSzXGUIM/l7tQBykkKIIeoAWUX3mQsOMQBz37KJNLx0QIa5OV
9cI0HO7qAP+d7hRD/5m/FBKj0hdamtuK5rLeBnayNuZbDofK79enUrA+Be3CW9424p8HP+bXGMoU
b/vn7mdNKffUcafLYpew9/+aFcubmDCmraJTMi0YX1nGz+IXWG5bzr/a9HKg8MNtPoc/6fTwc+tW
i0Q3CzQ8L5b/EztaWybRwpgRTcyCqtuHO4tlJ14ANKuEaiu6aChmirIHFvQ/QevrpQxXJjsWSjkJ
ESWR3hPJqWZsnlSn1fcsSIRuFafo4BBSvs/KQRPOL/dfga6CfsVoASeOSOjFi44QCMQl+8xABb5q
F9gi5xP4IK5tBoY2n5T6VBGFRbOFPP7DLLialHQLt5lqUYDzyGCLPjfhcn7YDbkkwyadnoGBCJTM
EfsmkpymGK1H6LdHgLAm3AwjcOPUdasYLs9q4c5f3fD67v4nffNrkFVOhnF2v89JzdJGyI8hRdcx
qP/XBN+EphXnf69+PuBH6sdAjpwT6Qyr6TiV9An99UxMu5qIrwvWCtUTxlCE+f6C1lfjw/YMT24N
cdDmwlp8WZLe3ov5erD9DpHHZlAoJUIOTi0vjk9rosw5q2+xBy+MNRSJFSKCsmjnf97HYUW30+w0
uFJpakYVkhfNtYBOP7m0teyU22vaGLiyZDCmqfRTMMn4FjEr/9G196st/sTywGeS4i4FCnXKVXWE
BQ5gflziGx+gy+3Ag3bmLhbozhq382bafVASG/uIsMh8Cw3VteScGBa3Ujy8/UPNjYtyy/2FTP6u
ol8BXEK9n4FKaWQuJMeDahh+rYfomd3e2CYYIoSVcwj6Hx+Jockm23N5+0oEHd5YJifvioKkO5s3
TgrfYw0blXolXHXTjrMbw2mov6m0CImCTH2MLoqhY7J5FfoxqucChHOg/fFKEVZK+NY8sgGm3Sle
L7EX9tkPT8Q+guWp2B3MtNDikaDqAu4FRHFiUzrBJQT3qzOz1isT/jhVTlK6zSlrmcpNpPwQySES
ntuslOxogVCGaYZCusTTFVEiyIvyNukXk6WpAr+aVrjHrWsyfe6TCp0/kd4OzDe6DqmYmAk4RMR/
SEsRI03F0ben82XbolACcSCKY8Mpq7GNxP6o5CjGcahYNDGfdSjscYYcc23dEsxca2p65eSGyjD/
S4D92b8RaXWvnoFkmi4K/FHaxQqTIte9l7p1rihP8aaGlrsmZPUDH19M+kfDAol3pQ80/1j2ptb4
E6dZ5ovMzGayrnl2bVzbME+pXZewK3Oao2PtdYh6LgYhBT1oEAqLzQo+BzYHYPqpGWuAwdR5sX94
Vbmllnlz5cRFN7kw7RDJhmAdyVvbajbfUox7ZBMmqzSjEe9yTLl96Wz2mkhgTtSz//4G5WMEcu52
nJUIq4EpdZEhAY7kVYSdeLBlCwAZ5eYrBsnna5HOVZgno7hdrtUwZEhN2PKtP9FecgVm2n4ckTo8
LUJYhZ9U9UGz+jm/CQXZuiWrjdv9g9yXioWWHfBon7LwOwQ2VolTWziy+/8cXKWCJH1UXTiC4BGN
lcrJKmBuYh6qzz+f63JPpdgOIHcinq+7V/v/BcTGboi5qKQf/2zhwsj86oor8ppDhFAVJ0U48STh
qCKVaGH7kQjFoyULjBZVAFX1xDHm9skqCOX1qblkfJGEtpnzZDzvIDpPOJR0AQkcKd/qeyx2d8O8
M6zhBdOD1efBss0BhC7smLaCwInbripyXyRmk1e1GGl+wEkCQnDdnUv0wRErFrhTPdzSi6442TCU
zShKZafRFBEcVhLzzbGQjk3MtlUA8Tw94kfjhJbGNvTPEx52gbpM9ZfsCOPBZ/Bk/T7fBBzkVJCK
k/lr7K8pem2FnReEI7bS6/ZXuQMdbyuw8y9X12OS+j880klg+MRQL4Elo12dqCytXzL0u2yOal2C
AR3hz0e1gpysjTBaryqV498LM3SKw0MPADZ4ejpP9uZJy8wAJ4FhmQhFkuLps9LlVr4f5Sgaw4n4
es1rd3wno698E55arblG+CmSNeO/TNzuoZMcvehIO3hIkOdYq8A8CM7k6HC/vCw8X6yf6M+wdG48
YzPTjc5hFig6q3JqZATWv2mX9KGSTFyaONd9o1CP5O7dJ1GcLQO7zsbL8hz2hFkaFA2+pTQS5rof
Rw+fb8dBaSRUMyrCOlCgjoiOXsycnEMtvKNXfmCCrm4Gp7lhJARGoh5QIYsR4Yno7kbpDfQQR2wE
fBUs5gFguNowhxkNVlCh/vLbw4P95Asrr2zKvp8EqFvazk4DWabr15XA2uCHw+iE2lVhyqWhSX3j
fHN/ycEgrewF9BMkVL1wNOLhqy29DqKdDc8A7xd+d2cS+Q1AaXFeCNzWxfrv0B6vJXGUvx0fgJDo
gJUZ63RtXRAQvK2zWOz0TaNpkSykHZOMBNneROiWQR7qIgtHKYAIEfKXPK5RWml+GIgEQVCAlHLt
0hbZFoIn5kQUffgHRojvwduvqHkt83YfYIstv5DlJMS/1nWtGqUvERFmFVMqUeVriOXazmFsTYwx
N3sCYZyZKhNGunDe+m/vFFcY5gIHvCWI68AuVfaRdRooykBhOjsyTTEMaqQE3urCyvB/IWUXsgo2
LFNMPF5vFUWvAfM8LUGyK9izJHjgfqsc6JlPbBaug8sdaEIEUvblEz4eO6z35bpR3E4ztA3PRbHe
OH/1Rr2+miy2Pb1mcVRCX9+p1PBvByE/7g3eycm11b7dT9RNM9fDXTmblLS2v+K4vwa5myHZYJ3v
yaD6fWdOCq8b+DTo5P4k0w9w4vrFxLzGo80ENlwTCwnWv+r1FNlgBsYThe2ZrKW31vDHQrdLAWKo
1dMASNq6sZAu+af+U2uXlZK9h/ZRsVBo0VvUV3O4MNW3zJz0Y9kMgl2Et6xUpOCtnFqP4Te8AX2G
xZgZu4joBSn9BlEIOWyFO2SSPbO4Uu8kQ9Ajn8xg5NQ0Ge3GsmiTmd/yQOHCEitx+EqqxdY4ceDA
g2mkcvWJXpNGePl3lNIdLvS01u1w/rwFgCnOPcxQHCtPAViEgEWdPj0Nb2MdyS6T9mssM8xtPqsJ
KlpGb2UsprVnTuwG1lJUKBZ+AMb7BHsANMB6uUkIFxK3PuiQpLWRedIw+sDt/BZHYHVIZFw6UY4O
KFUYbH+HB+X/qwlJB2u4m46QnTgg+wNeXqLNJFEnQTF3pHpXyL5BJOHzEDYM5cblidgBLmnBidH8
stPj9Qfyg+Uxl+mkNckPnGhzShKSrofWvXa5T9Elxm0H8CbAH7Z2WzLnElWDRmb9C12q4gmXCp18
YPliar69VGhKCYNKGeV1AUoZqQHJrZt7KJ9UsJNt7soOSy8XTv4ZiLwW1fkCb4ocZV7D87dGNXZB
hw+yX6JKONRXfUGFwi4RBl+96vBc3TjdMGYqH6jIi+aqDkntF1ffzdPfFWILoZF+UWhZGu6t6Z/n
CiT3lXXMTX0gbIgg94STa0ZfArAIHUKoiozN89CoU+rtYf6mNzYUW5gB3ZkGVPYhU4H2IGVdcaq0
CT9u4V2uMREw44Z2piBensF0FN5iNfIJy0UmVti1+XvY32BOj5FHqhgdFLPV97YnETVfu+d3Aa55
7ty51xcI8T26p4ZjmQOqBiHH4gor2dDuEHj2L/rgw4bchZy5kQpHXZAJwcdudXOV5ruShvJYM82N
3Y/uGpB00TbUQKJ4cBVjbHOoBjUrT++MQGVrj6B8sxbus7ox1+e4kXPqXle6ZEhmXOL9PszVPdtG
hweRgBsHWjeU1U4M9Mud/JLMd8sTcO7Etj7pmghR4mmzvIqRRDKxDKiIppHywSG8FErVEyilggIL
ldHoWmnuqLsOY/JZZah+doxHpmoYQK0ri2n2S/1cO42d1x70HQ05HpMzlQi2tFfBD9xcnNB+ekLg
Yu+v9mmu60QSYvsBt+QUhCjpoPNZ2RBOsLZYaqrz6uOn49RaD1ib1dQHZUdp3pspzD/IZOt3M2+F
0uyMzibeGJPp0pT8kRxS4H/RAn2NY4TqJPmsGGs7Qmh1kYK0z6tvgKWUs8ojF9LbuJJi2k1qH10V
i6cqpJwfE6Al7hB3DWryREH2ynY+E1uTCcexbElgfxANpr86IRfKxL487s6yZYk/KFoLZ8OOUiy7
c38nVk0J400+6rlXD+MGEBRvRTboPsAHcMUSWrayNc9ZHUZ/UnXDRIu38YKzlYxvsSOqFufLLoW1
4tslUfGHARIu57fDq0Ghtv0spnWc6MS09tVi7evAWhedshEMLLv7T3mq1Xw6mjb30Kr6FUsbcX8+
gHgV69CCSnCctD/nnWqu7YVnwu9MMvVguFlpxIxoQ2NC5jSVE3Qz1xsMVX5xnWPlkG6NQd4nzSLq
hgbBypE7h3xBreVRzNCt5tuaWcrE7lBjGOXyW1KVV08/A1hpO+efHKJL2bIkC8UXzFGyn/udOVVA
wImZ61M1ngPK+fgJ+pQEOL9B4tXSQpu1SqhWhllR8P3Lxq1EDwN6Ew/jGVMYNTqz4eN33BdNTB1C
wBQRAwN1LU6LvG1buwWGjn8f+pL0vrkXKpdjVQHFQnqdWQpDrkaOdGW76w1ODWz5GZtumBMYWW+J
gUC7HQObTOUgnGdQZDcBc+m7Pbe7NCroleO8y+q0ZupZ1hYerQbXFJrJZcLUoawwn2Tbf8XUm6f6
SDX9RXl6PFy175koai1q7ViA8cG8EzTSHWP8AXlwVNhQfIp/05AzgJUqc+W1bVSSugpeVY8oTagz
PdSw7ZgAN9PynD7Llexb9zIzYuDEqJeforV3g+fDtQ/rb/wvy3jxfx+++bt724ETvsrVW0t6UFQS
paAnZ0p9/fRVDMWicaiDaPXK2SoUnDuZPwUo42ZbDhoNhSmxPmWnlH4P6rwDUPHY+a7IP+6W+7co
fpSaTnWEW0Khv4eXsC1tDu777QjuhtesHIo5aLKyIOj/NOgpNNWydrtwSdOb5W6Aj+LkadvtacCb
nhsoe/0dEtA6BtMM7WWM6ujddKRTZx8HJHhw71+GdZuJ+U29jM+IsPauqT5ig1AoHx9kmvGuviqc
R/T09G2xlgHUG84hFr8RRdOXE95tV00laVTRYts4qjpqyJV/eQS72Gc2p8cyv5WljLG1oq3Y5ItC
BHHGp88cOGz28OKx/omEQxzFr+SwjJDwvManEJPNN0tNfXzb9s0PlgG8gYi/bV8jKvhhp91uPayr
RVg6p/kSU+foLkMl3Di2s9UMVJ8byIDNen5Uc5mqJZlC7t4fG/PM7FC2s+v5Ps4k2VSwOGVquc7k
9qvzczRdupJuf5WabD1LPVcnWIxeRu/aJy8mZBPx6gKKCWnXAURFVbilVgg8AIdhpp7UlYDPArgF
Lxiv8Nt3QAxZFE/4xPtcElwcL2jV/j4YXU3B195miWUvPaDIji8NRFoIfkpXTEoF/HiT0rK3VUiz
AK9bRPUDdBVdyd2HLqsMNFb36sMd5jQlcYbyffSBeLoovfAzP1K2phtRtTU13Thn+SQxXRNrN3ej
C/jjOakx3EweWndOREhpcIETPXTgrgpUyfPzMBS1O1d92X3q+orJkm4K6Tah7unxMP3eGlZdPRL/
wON1AJmWjy2lqa9DQc/eJfh8XwKR/PFapZ4oHLkWsSgCYZxlzQptcBOi38Jnyq1Y6CV+vUV6U04H
Vl+Ws8Hs/X7nor6WcreyiaV9es6KPUSgXkojyo2MP25BH3ktKYEugBIS0PVLnmduIzjFQiIbdtl4
uSSLVTo5AIVHS3ycnstSM5+fA1C1IY681mpAp/m4PzKPQfg+z3OMTi/01OLnzXsL0lIoRQkakEYJ
4CMsBMm6egs6gmDJJOgUB08gDjehIiRz8fd0TWyZrPOmgyd2CoVjL4VRvwaSmDaxhB3DffWu8teV
NPSUgbQYlVXzTXM0iWcx3/OF30PIYD6f28fe0UZ4FbQpE1jNPIcUvpgmFRmciKf1WWI8tglOjKTe
CdN5cBn3L0qVuT/X74rt1R8QE4Blk6sz14t/g5SbgIaURsOCv1eSremDjoNGqZxUGqPg2f56f37f
O6nUKJEpfF8y3T73csiGDpswkI03fRyZcmHrWRbewKE9f6TjXCLsO+N99n1eqNErcckT889ApX0e
Cpz6m7oQsw2TZMYy4w80nrddVurLiXE8tIMBKUcmGQPVuNLF4jCmawPfXxHTmdN5AjQGKclczMhm
qVbm/Mu/98ipzZLbYGx7upJ8K2UQ1LBObjRXrYqbx12YWOvJLVp4CFR+CdUtDmgpnIgmf1gK6YUX
3EIg5SP33vcwUc4vO1XBUooXGk0j1ZUi9YWq6VJGQAFsT1Hvy5Elxbc7JX7rt2lbOxToTesIXLcv
D+EYzE8XGKTHfqNhHmMz/cEm1REEcXkofsD5dMt4viWteFBD9pE4W6NXX3RFkRUKALUd77NuinHZ
ggaUyyq3hGHLAj76yVTGvOmjew1uJyISywdQlpWGkQAfUbfb+XjTL6P4f9HFikC4gIKp4e0NJcIE
9Vlrgd3VYJfRpY201I8LkyqKtw/0s4vk6Qv+GyHKcodM620FjRBnr+VDGSTSAF9WfU+AXkna5Sbf
g3lf5WIJsU4ogLqy98DuDYFJcoS5t2Xdm/man1YSPHcwRsWPWB3YUsUEM+DW4PQGNz3z55Qt69Dz
Ckhf/Wl32e72QX9n8tF/Js47LvGP8JiTDBb2/RRCpLfXo98vS7w9jwtuW2Mwc2WXJofCaMykwkiu
jFJDopQF2pCayKPM9hHR+P0UcpU+2lLCpsv9zws/QhJTTnKyS0nZEnGsntyWz5ZnZpZx4f66ZK7L
0hP9e/TcgNIEIFDDNJh9Ke35/PNSoe4TgNSCvJ3UpYpU1KcIY4kgqiztPxnFWSS1tyl1EZrCv6eM
QaKewfMTzokGkrqxJ9+DxwsIB1widLgzEWiDa6LNSCgbwDIBpH/cjzUp3XxOpS2QO8kreWLwWd2z
69ds9YWDvw9sJ8mAjNwRTKXl4dt+Y7jKWs4jJuuCSopV/3Ev16i9540LBAU4Wl2UIBqlqWw+8QDT
x2JxjT8Rh5Cq8vx77jxsD2OEZ9zkRtnur3hMWXeTfpJQXdcZFrgNdTndCLSq/S8UYTrUqe4g5MfF
iNO7vIaMil76DciltnS3OC0Ki7jowZVycHELKQzFoEPqFsktFtTrfE9H64+ePBCoEx4cxgDON5ou
wH5JcdBtJgrQCkUqMhYflNjrY/hd8LmUEDt86u4pFXHEk7uhZwrpBC7YEEtbQlMnku2h1aPyaLyX
5Y8jO+baJrrAhWHn6LmSB1VS2o5cpQDmyyg/WUPto+vJw02WoRTbWxZrRkCHlObIaNwWFjffP9Nv
pCXzQ0hk8Hg55TaWCBO5dDhp3gG+pZ0psnPgKcOMoBaakadhXMg72HViFr6j9nyOnuRTb2BEABfF
tS0JpfF/JukQIxox3D2KHwnGN6CE++P8RPtT2Ku6pAkStE+GsdCzaT2mpalZsNjEQQXlB7K/npnt
iWurEgKoYwkI69rszfZlljAiIyAy926hbDvYT1KOtlfpPKGyoHOAYcy7yVmjV5eVMSQ0ocewdcUc
zd9QWmid3ikPGjPQuicPAPDgq9HoZxnRucZrtCBZhAK0udrRy8eeJ7c6fOmctexKAlkh6YUo/Yy7
3dU1DGDZxRaEH9gf1/f8hBtbOJOfkZaK6RHPlYTsHrYeZFjYF2zBJ1ikdYHoc5CDON/rz5LrnU0T
HJE612cfzJc2hJmnXN/6bya7NyUJ+oDln2JEUz7YH+5sSgFnhs5Sgm1l4kDjkqFhQufIqku8hDhV
on3o+9KCegfai3RYwqR8m33Q0PHOPb6zWYoQqCQZ8CgjunI/1xq866Zq7Ao/sa51ecZRHIKnIAww
T4ZFbCOPbVR1A5pCa8iqfjM2C3+tQnYBm0L6AloKecrVnUHUzlWaiZelevW91U/H6e1EOY+oTdsf
vUWvsQV42lW7rf+g6tCRWY7JbPt0PCmLS2ucG3tpxt5b0cTCyUymOd5jCQjBLgnROBYw2X1A87YZ
0imyRb8i75iqJedUGFp2VebAm1AdUkNZ/dzRcXqf9qEajIgoPGwVzgMDw4Eq0nf9NOyI8l3Dc+Lh
WyVLWTwk02ZjY5mDrkOCR59zmIq+Npg4OB4k4uK6OEmihZ2QCDIm+3wyocZRt8h2SGEa2Zox7Oon
U00w62h4uKC2Air2lHYNd6LGD1jqkoEgtqu/3R+CW4PLnWrRZDpihfjkYmWSB74P4eSceLEvwnTc
9YUJ2On+TxMdYBFmdNYdg3vZBL5FUNNigN6m5lBXzhRuYZvGTRuKR2m6RXnhVoOOx/yYw1UqWXgN
Apkex34sWaMyutf1U74S6lF6uINKJ0XoKw7WiaVN6bRTEd+nIf6bNpUkY/EmTfPXKDERj8uCVAgI
8Flc01ztulp1a/FRthyZcMiO69OOipD3b9qlpKtT4ddPFH3f2rmOyTEQo2OVUO3O9Zdsl3T2cH9K
XCi68FLd/venk5yDLZHA5U2UGhMPewaosBam5ztL5MKaD6N37+CyAIk5I9O4mJ/mtdyxau5pFacx
dJPR0zzZIuFPP6umWYkm4NQGnERXBIJ09HUakAA35sIX3zWQ99lVdbWyHf8aXjTZgy5OUJXXSHBD
YrfPf4k7n9rn6CfhHXPreIniv75drCUQM1fi0j7ATQmvfM3Cmx5cTm1OHTfDRe5H+at6fZW9zqAJ
6TZIG5jKMaIv92HK369pnLgcSqjc7gaV2697CFqnpYsccA+qq34PSJMl2qSajWrY229D+mBo9Wcg
MIq4KXNqSMcYrJ8gLOp9Nxj2jKg/eRJn4QsnXo46+ZaXSMpAaX720HUb2IMO9FJe7/PJfygL+UhB
Rt/ZWcRsMvnWDN3IABgdvV/zOKUlq529L5uPrf9SmIgpO7KJlaIB3PlLfcXNhBgaR/jKWLcN26Lu
EbEhX82i5vjHk8aA+ALb7Z72mYakib0Rj+geBuJTTMdoMLrzNUWpn5rnNqXXUZbWwcwDtSLe9Ize
WtgMFA6FG3jlZkwjxb9ruuApyuyhXiIrKojDAEtjVVTSVGJAPalqX7Oj26xrHKJzxxeVMCjTlqH7
GJI01ldD4pyB4K7vHF6vSx7adWWmsmwSS2K0fhDe4SedOXkmxd12g+BkeFGzVaA4SejHk9eT6I1t
oHOlWArYv8hNA2AX4nwuNvrPU6R3snQdM8KPU3bNU5wBB1e9zNA3P4G+N09j1eXhaY66XwR8Kqj7
SDSnFzf/l6xhrj/xAp3pyhzrtHusJVsXCRffYDihwLaQ95MqrDoUPy16c/Nd5o0m4hS50eqC5Bv2
6WOGi1V2Jpbjo6VkR5scNfjWVunVr8wjpX2PgauZsrDBJBZZIhp3LTBiyQ+x2V1K9ZnvssRkt3zx
SLN4Y41HJU79iKqDVQaFxAVrJlIYvRXqpHfy3/DejsFRnN3TwoH8ouc/F2WAHCw6RURHKOs3n5OU
QwGCpuqYXWCGiGb2y+Lvpe6pFv1eYDpCauh0FdTYrfD/YshqM2WTAkQOJnwjSiGiD9ifRID/R978
0G8j8GQKaImz03xOSk3GJfxv4AimU/UPtw/U+EOXDZvTVx8He88mq89/sdhzruIfWggnuo3fW+Ij
K6ildNrYAuui3GtoPDEKq0Cu+bBTtVo/p88VpKY93w9ar9mxJOvDKBb6pTnP85B8TaKxOLAVf8Jr
dDiqh/w2sjely+u1rxE+qsWeCIBg3yQhxBl8DHdEdafDwwxaM9JGowNmc0w00T6Qu3NqI9+XQGXX
IaBATfXUhpHLA7FQ5na4eevNIBZz0+yCAgG1NDWTBQHPVoDYwyb5JrHe7LHeFAywK6t3Bb8ycf5/
ExKuMScB3ls2BjWopYRbWRzmb1LInnlMt/1bZd/2A3nBHXZm+ZRefDxdDcp2U7MNfeh9iQwFJaLS
ESYkWTqS/iwoGWlB2wNuChlNItunroRp2lQyMl2Sn6CmEk5OkAXyEpB+cmMg1onutEadaOWltuAN
HXIbwyvYFOc74hN9S6VVqRK2Zlwe+hDfG4snS23JRk/DglMScMyNLyylus3dRWO0oM98X/k/PTCI
zRwGHBcFj8o0dvMbnlORrDHQ8u7Y6QrjgYOne2vzcYKe8SdxBnfKxSvQ7PSB8nnBZ8JZ8+sGIpe5
Yh92oTjNEZvthd5OaUSOf/wpYVz7u9OuPCJGyoC/PYYpsSi91b8gG82ZGqvC1YJ/L27+0DiVeuH0
X//gdqIsaLpxvIRr7B6pMP8cHPSjZA/BBFEPsDrDNBOxyMX8q+E5xG31ElP1YSLI6WTpKzoXvE2p
uBX5hEFF3Z15jWg7vD+cwUr0pqs3WAFHRhqCzyA6Hz/5AXd/HvYKK/+7MDhQUo4khKJUZxjU8yz4
rjHnws14eQ66CHsk4YXvtKMNgJT1s0sR+6p7CHSQSfg47Cjc0/MzMPbmtkNhP5G5R73oL/hZ2T35
BBXqlw81K5maZk6x7gyinWjPJHefKoGtjfPew4R/x3rdYdvDkXOzzznnl+7pSAoLHSZNlPlTPSpC
4q6TcLOW3MiCEeBN5epzeVpJIKAE09pd68QuwKttHneQJrLVtzS6pcYETE8XnkgT7ZaxSL9VTPmM
aUgXkSJ7BMebCPseF52NIWd1YsiSHDx8F5HknWJZ0T3moI/PesG19sgm9c+wWv4ssMFp+dJrHdcq
xSAFI+Ri2ks6m4evGtomX1CHQYupxq/sbBS5hlqhNElr6AZw2MyEl+rY+e2/KPwh1P12YgWldooS
7YI9ERa1XTq4rZaOyrZX9+YfI+IB+a8azL40hQGAd+w14BUpuJ6YssF4XmeygUYSnBWvjFlK+Bjh
5NIpa1Jfb2alf+H/XJU0oOzBcqwbpSwpFvuQAtNWejl6ektdxZTOfblOoPDfNDm14AOmJgaDyNtn
gh6YOttGzAm8gQx065E1XUdF9NXu7rqtbqCrkCk6pWMymlMvcX8dM8jQaZBRbtbxLaGUsG0kimEk
OlZNk+cEaIqsQ7ePMU5Kp5DvzYAhc6yiOgFVqjYY3kRg3zu1Ji+ZKdjJHh9zfSv/4dFwScmjf4LS
zoB3BdwipnvapSqp+uiYiLijUWZ9F3K7ppdDGema8sqrlhLKF6NqwyJEK8tnL7+CjFZm82apA+RM
1jQqmLqjmShMfgbfOpicFnJxMxx9CjjZhW01MfRfs6+LRuOGdxi1qPQYYYwbNEBnx76RL7Tg+3HJ
dvPHqmenPhf7T8v+eS0yfWMnsdsfu7+ZyN5bw0CRIQ0xJA7Di4WaEy1A1rzbHW+e2KsOth+gjy6r
9T6ZMagerefu0mxRV2vBsW4xDnY20ZYmkBPloigmezeAzY4jVQUe+6UdNjKenkBQD2tiwk3GaRrv
rcl6JwRwEPwGpNJ7z1mtfepJW/bBBtSU4jKcg06hjTY1aHF6CpcnNQCO7LEkEKDUNI4nIklIPhqj
hR/tClz4yXqh7Jh/2E7QJWA3vfBA31ptiZiALxIwgVFj3PFIEPS5mzkJAwuCvCc8LYzZo4qJ0Aig
uavYejTt35RpiPmnvj8iR1dshIXhNkk7GogaRSyIbtS4O8z1VRq+eshC8D7fc4dCzb/udRD6unc0
8IfARqN5hyAzQL8RvXVDTyAIVZ0uFkV6Esz//B/dR9Pg9Z8WyoAg8/6ceScAJHnJ49qkjw2AlLOR
2g3oPeDuJ8KuaVCaHJDZ5IaS21T/akFw0V/Z8vq4UsAG405aClc/+vBDC7Wx7QgYjkHIrcJdW35l
Ai8AQYKzMI13Gts2fQjsypQnS0YOyV8ZFq0l7LcFoHujU/q3rZTBCrpmpmqc9fIT4rltxL74axLb
H/XVetuUVcP0J8NDdNQeF5OkN2gUy959xp9cOO7tRewnQHr0mD1UpRSCNasco6AwKyBd0qeUvZ04
MaIRHu8hGQYt/i7P3YsxYxF5+MUfWp+YKTtm3doRzVo6vdn2hzKCtCH5DfKbKxCe37ohgmwzf1rz
3RkuO0EiIYjt4Ra6iCUxgRhdtdjrUbevtYAMr8R+cAuM/FdNxsMvZQlM1/Ksk4f39rPi4HPI0JuC
t1U2ny/iOf1a8xjVoxLkjiX5u0TMEEAWl1gbNGuo+yO6CEPESKUqP68x2DCsI7gHVmVCjPT2laZL
619yBMRyEtKQiptWHMwy51yPX1JjupXiyL7LlCuuAZUtOroYeIYltiKwWPuF2QQqhyH6g0E3U6A9
LPKnWHp+21UjQP5eeEVEJYGmzY7wiopDKfPSZLHm/ei23DQIRazH9t3kb8fhTMzKxjXx5kvLlnMK
K3GwDWfu51TSbydHTTvK0yAax7/6OIbvl6mxOjjEhGL22VJAJO8LQ7syvvea36VCgwCTXVOx6nvZ
mvxPhsWwgNKKk8c7yuGak7vnV2dCL1wqHa6qKI5vBVoDvF5T5vWPgt5zx0n1siEnXaGL5Ka1vcKJ
ej6crWBC0wLZOl8oH9SNDiRizIfM8Z+HNBERo7Np26rKCWBnMamaGlw3pnx8ESk/bMtf1zRYuxVC
A8BVTwRCrcqg5wg62X4xgpDbwLeLCiNITnHjF1kD063M1OpAZ4p8CXQxcvSwIULg/aJ+pbR8bLOj
UG47XObH4yjW3nJr1QpCds1LRSjkQFk9lWOnAPNr9VD+55gdLZQML5vlEVI5Z10118zH58GreP/i
wuTadvJQVE+L9db8th4Iq3kBJ872frYzSZItDnvzFkg+d4UqhizS73Bckcm3xds5JbJCuMMwfF8Q
v1Rr/z7SeB0/kqdLzsyqFm3Ohrx/bTVovRblhzvpSdLa6bEKAAltmPgEeUNopoDbDxsCutAXUq+5
yklPmvwj4NyYzB6Mj3FUYFCndqEYhGZzZGyHVo9XsSfeUeOYiqAJ8fSe30bVDk5NUaMoUL6KAmgg
GftJ7AYyC2yy6UdEnlerNzqkIQ76BrvRllov9TfUlUGxhjf/H1sQ7WPrHLpLDfrqJJYV1Ro2Zqdf
LXtRB8rN3vzMt1tXEmBoNYOfa3PXOMiNvsate24K5NKO+HEC+vezx3PoNIoeeBlU10emnk2RUT+L
TBocWWnUUt4cwCaylilrBgWltwe5eAM59BN36YcSbeCtSgQkMml63/QrC/AAdYVDN2YhnDDU4BIF
xyI1aN7aJhP7gv0kDyyVRxFy06rVuQYVMoaUD2fuS7RdnbaKhSIcWJ/rb4O3xBmyQdna0Wm0GKtw
w3I6S8rDem5mmvIRb5ICwtF5DR50PFu2z/2yENW/5me0Q0c7sgjDtE10aTQfm7iaXtyVSizsHaBg
gBPGN5NOe2ZFqw+RsJiF2r8QvRSQbbRZP0T+ft1S1OBkcbcLahFYPq1sV4PAeH0NOc/HAEecU5Pu
1jbbNCGvmBdyUg80CjaX2HtrMmnPzRQg6GSsgD/ATkf62TdwB4ezBodKHhMQcrrDwYi7fExUTwVh
T/Ffn+f2nskVKg+P+mTuBkaWIxVG3P+CQ/RuFYE600kQmHLhul0Fv+hXy5e+D5M+77KVv7mPVVCH
4gMprye8qSk979NyLJXOHix998MQMdEW4xFreChw24M5HlgR37GDvZxCTehiTlJ5PV3t7UBp/CaX
fRVMJ+nx3qpWqSlmFomdnAF2XURhHkhaUR6R1l+mBPYPcSeuBEpZK1xYB13foLutAPVLqn8iPHRK
pC1PUdbSXYRt4Vy9XPlzq7CGW7HBNl38X1WszIP8m4Fzszx0aHe2QrM8xs2EPnnbCwJWEPnaUcVu
0hqyKFb2HCv67GWRphaGQeGUtgNq5TAtEd6I0y3Y+oLP0sDfV2UzPui9I1Q0RhRgiy6tpjKh5dxX
yqVWOLbf2zUdbhA2Trja/6WA2kUz/GN81K1wTA8bf31Glss/cuSqnNXE7opO73iy3zwQwr/jVUAN
UH4+srpCT0tl+xHb6aPNvTH6/8STnabR2hP0b7uGxbmMquKw2aqN5dukwzDKvbyOBEZgmBGP4+Ul
bA8Rpq+2WzIUoH8SCSuHv2pTBcIKv3ovAgimnyfCBMNZ7bgsj6WlBvbJ34lm+hY1JWRjN1AHLUrv
7Fmd9DssL76jyQc/eLwMs1Pd8KFr3k6zY3QGdMprJFNcVUQqBry9+E0GhWFq/z+mvWuTGk7eTDW4
6KVRL4u/Bw2xRMy+qljQWc6Cf2yYF6K+xbcBAhh8vOeplSQWlK3CxSK0IJBz2O41Xu0B8v2dlKRV
U2FFvR+npRbL7LJhtidQc0i3yMgjXCJO6RK1oNnV1NbpasUsJHtmZSX0WiiDPYF7o5N2uQ78QNfG
WY2jHaH9iJ+brTuNpmrwM4pbsfEHCbgTLlRw3+OdTZpICDyda4QFjVDSL/8u6r9gkcxqqjj0MiT+
VeznPiShiKPE1s5tiXObqOClpo0RZYDSx/Rx3S8jIpBr+MwKdyIL/DQoIY7F56EB9CIG/UdlNZ4+
mCXjeEbbNrCm44uefZj7Mgrnfc22/qYNYZvjq0fXT/dhSI+oYQ36eAV5FMdr3jLYYN/taxPW3w7W
J37w9zuE+KqdzSpvy46DlNhiUl2E3DNGT8eJMZMWAtz3M7+2CiYtpShy390Ibt+ko6iS152DLkur
/+hvYof3iY21kHDp/R5eoH2lZrCUe7kKm3sUy+kay474zFS+HBH+o7wKnQaUGykumSykjiYXwe6/
M/VkD+F6udONv+tSBa//2h6ksmiDwVPIgbujRWb42mLNZDj+gjZHrLqeJyw5F5HbKth0GCPXfYmp
zUpmNcJ+ZURGCw1OmmCKS3zhBI4Kojwp3HXZy5WqfEvZBRFdxM4ze7yNi2I8KZSW7w/uUn291VGw
kL7QjEePVqhK/twceg4XuIbYap9++ZdbUOMSarvgS9Tq+CxQr0HLqHgPVyN0o4gpqE5F0w6j44+Q
MRTcms0fStt8Glg5ctI6Vf7IGC8nmJ5TWyCqKlqMIWEF/kzyqtQKAFTZIi8apeJhsavlTlmNYped
4yCU9mnu1lLkLi2DKvs5NDd7dJ6KEbi49WrBu6YR8yuWAh2ZsQGbVLntyFQG+BKSLTEOUPMJ2KMW
0e3CAl8Zq1TvoHZ3XOP2hFzxYWXsSkdr1gwB+iemLL1z/YiOSs0LNL6k2LsI1ZiEEaoetIiEaMiT
SRmKP5cRgoGPlrwdhSuBOWePDY4E1C2nEdJ0TdtXgM6jfp8NtyQZx9ZzA7weFo9HVkFfY+r1aYtG
kULiD3njHd3vbqkkexeXe26vFCsaPRsTTodUthOcTewJnSBfgQRojmxHQSSKKVoTc/d0X1/kB6eb
IyqhIk9o1xk3nNBe6FN9BJl8Yu6MIv/UnD25kYDmsrjcOIbyt0uuM7fRlFq9HGtMCLVXzr/ylHbd
NanrdH0ZG/vUT8WL6zqfYLsYmT+Isn9/CIm6/YRC7Zx4hpDWOnJqsjxFQyNy8jQwjxcC6L8BS64Z
72flsCw5xg1Gfdt5CN+fPYhilDiOxBc44GL7i2gvEq1me4wFYBNmfFoOcBz2JwYdMRHtpLD4JIwA
uQh/J3oWSYanrsBJA97AnJxHKDTmGg+25EubH1ll/Ag384BnycFJnFeTNOyX6aR6ZXZdbjNyz0wS
j60Uhjk8BIkwQY40AkBDXpBN8L00gOFk7CSIk2Sru9tPOOWAKMhGsFM6bapRycxrcaWNRgHdP6En
/IfaeE6XUfizBKdhsG5/KSx4BeUTS05vA6mZYaTHZhiSRv2xbRVfyu9UfrNeIwtpaGM0IRx+15Dh
4Bad5koryvIZxvizx5SALA1fpbwMhFYncE7HSkIUKI4oUHX4LQRMZeZpcEgcVVudCllnRiNdyUXv
fuevXpSZkJeefm/2W12K8t1qeYxsBnf16AIsCZTL1XGoCJBRRv+NB9bU3SoPQNpIIcK2pk89rQux
PYbl5xHtpGo/Ejbc8u4DJhvHrfukxfAfzqPtbzWvxtyu6ZC+K/qeGNw1GrJ2y+boox6qH5N8u0xO
fj4JxhGXWK3yxJuKOXjGhd82ewtX8YqorZZFJ5ep65fkops5oV/xaC0jfdAX1HNxwNwQfjbztwZn
CV8RumFI4gR9D35jNIoaEiSIl/zOYrjOmIZKURMW8UVcSYP3wx7+46x5BqAPs734SmzVSJ8gwfxd
FaQf93zKHmO57aRLI1BOoKupGQ69kWIUPc1nTnKyEb+qNTXSjyz8Glriro0ZGrHMs7LgY5etbhsf
dnB+TohbKX9WvwB+GkKqVDf626sptV2yTNaex3DOLuHRitCkErq3hIJGCvzYz8JdHR5ms5ysfNPU
K3b3jo1d280xM/m0Q9G4ln42Y3FEvkgMLwfRIzF53naKYRGMOGbWfoN55oIDsUvz4AJKkzIAvU3K
GCA4QoGNSFrfcVkddLp4q/wR888s6lGHyxh6HuX8sW70K7Fyqbz/TTUBaNhAh2iSoYvhI1a8T81S
VoK4S66NL57ec9ZMn9zNeVvhuex8cq+Kyh/AXrBSqwYnVljCd+yo1e47PdvpYkeKPAED8RKABr0Z
RPjVVXx47Z4tDaNxNS39fRBBRgdi5kaplEnHl1jgTtpyyvNvLzNSljVZrHV0yei4B4/uU5dM+bS1
+RT3OBb4jHcJtassjL4N1AeYx14Wh+ERppn1s6zc2yjQfZhisvPXRl7H0JIcF/1g6HaxndfQ4b9u
9CQXQN1v9WTKe4FuvCeHLTULLhyIpaQnqGaA3WRepVpmenVHgRV+i4X0YD20rzQ3ZnDa5vnSobC6
TKKasw03aP6m1y4ibFZNVKgzI3SSvhIPBFsrz4NWejdfV8sDrxI1hFvb40Pl6AEvw/6MZ+c0gjdl
0QbhcFkTdzjWKOmp6ZCt/GrL2X4qRZyQAYlUbd9mnO8vviOc9dyh8jrpx6bdGhs7JB52g3K3dYTQ
Lhf8XHV8awat8pMhyEk4SuOP/NiNHCvMAJZOKde3ZIjFj3CNe+bE5J2gckQb0MlHVDy1wV5GF52d
rKq2UxkS018T64IkZDyHBItLoxZ2eAIbW2E1JWjZknLtb7eC5B/QVhJIq77YE99tnJWd1qC1l/kU
dB/n/kXknBYeNeJzpXUrMxq/dUfO/PsEvQjzedoqE3S9djEuuqfjupcaKivk44eBOQP3I9X39qc8
fllmASIHXPuUE5PqNLBzrCU5NaXj+sBqeH0zpjiu54oTZHQOV6kLqaqbL9OmQAyHHJ0SSgKwni2B
XVmVckhbI4sxuPZS+IogF9hOMhtm6Twq+/Jtvi3OhUJKRE3AYz2XZHnFkuYw/NjlhfsSiBybFirJ
+ZRgp1IMR2bBXiI3s3R8boTyY/IFtcanwN/qrCRSj4eaDJaUINmvZqSbto/L+EqQfItd3wTYPPj1
tx16C/ePBMKwrhiuU/Oi7Y6Gh5AoFWjIBE9XJ74VGjrvK8ctpQt5fCHXsp48R9GG6St+pyYM/6RP
2rYFevDf3J0qG5C+gHhsTw+Z0rwWsDNTDKzyaR3Aw/dL/4UaBARrS2y2czfOJbDPX1CWGGlzMaqT
rHyBGoWR7v6xX5nt6YrUo4X8QesXQWV52NBT8GpVzE1LtcWEVQcFWvo6TzaQ8bebMkB+lbdeYzYn
Y2it4oVBbeWkSzG3ihvbRotjwT/E235IHh9SuFyhX/JdT+TzdelNskrdO640TtfIlp65sAcveLCc
lOX7RoRVJrJLCxNdHEaDmhLYzqz/qJ3nT4aLwTWAph3bqxJsNLkk1ziejkzXRdRsf6OIEYQqYLqZ
v8cvei+aecKQRIgHf5bXRwGxIq+fEIHOswThVSYKs2xVWZz2C7SnYqriDoqnRJRlqXNfaKzOCsOB
1rdzLbx5F7zXyJD3m5BKAKBbjioiJJ8ydliNpu2KmoaOvGKS4I32IEWDpyUCZkWa1armsh7YJQc9
VDMNPTi8eytZUZIPYQjrvhw0u2WS5bEKt2Rdc/u7iue0nSofldwWQ8pzbT4DgLLlKw62vqKN7Srn
3jlxCpTcdRO6suBEubg0NOhKaLh+gGBFjnuWqVnC8TzVKDXWGEDBBby7ZWqV440MHvt46XjhDjuI
WscFHs5R9/C+sdHP2GKN0mW9I8EXp5K8aJaS8fyn/ZaAOFNrD51hkXkUdU7WvyHW35Gnj9zPuoyX
mNGNx81Jng0iG7/nAXKw9nRIRs3BCbPc5Wm6DaYcX8NLhVb9kjTxAQe/RV/P50TD4CZlXEadGODQ
vb4CNQL7c9D4l6WVzPngcxkIjw8fzNY/DUhCfvW5s44QnDceNIjul1JY5nbxqvDa2SO0z/Xsv+Bg
Ecv87na6H1X8cxV5oABFubvHwL/+p5BwBwCs0v3vV0Awf63RGkRarRc2M+rttoYTsl27oA5Fvmmw
8m1LnHF7hrPHazkkLLwHac6tb2tjsvBb6H+aUEwkfyDr52hyn8fTbU+go6avdeWISN2KcmfIeyCi
5HnhJk1xpzJI+sHi8GhDcfPJa+qTOiJ/qWtwX8wGmt8eMvij8ylEzZMr0n0INYI9TKKNaqtbQLV1
hnapW/Sz+HblkLZHZ21oWZK1VjcNJ3vNR8731urW2T2T2hI2eoeGvon1I9LuGd52aOGHxV+Vc7+V
hRDssQC52efDhz9pXBXLcGT8mXxj2UFQIYUUFsu0d4TdkRn+De1ArQJCiTCXYNfOftNPGUXrYE+y
u7yjdem/teNKSewYpSCnr/H5ztAYk2rY+ktrme6cXlFRRG1JqX5YBM6lS/iF8I4BJh4eki2GwyGF
PmaZwi96vZlEVhj4fOGTF+F9MDoTEiJJ1+eETGAmcLvIub14zw7zotDqh67dhg6SLrrYj56oEKwY
D6dbUH39HtjXf9w7YjzQZIZ8nE0WaYUux8FlIZwO7/rVQChq0PCe+Z0IglG3EogwPGZnAG10H/GF
duTACv5BnApe6nNjykC0IS/qOSZA7hxRtFcd8VJVDU2+7GyUq4pkhpmZA93nh2Bo4wlMavg1jpBM
3F+Lkbsgbcs7MkbieVKL0BW0ZCfV7pHmDq5x3ZPDXAXWuXkVXU4sfbyq3HCBZAAfHlxbEtZ7MLDN
RoIGIIsWJ8XUAZYo0w+a+RC+MzJIk1WeyPcY8WA8EC7SFsqG5C4Y6jr7bCK+KM+njHDLgog8zDzq
8E4LrXYvDQvrjLowFAdFaMK2apyTL+1Tbwu5AV3DcsAakwRjk4J1Ph3eCEm/X+/lYRB58Khq8VtM
NHfkuVEbLz4iTr2asFIuXgSp7VtFnhS1BS+Ly0ZLBVYKSfgNMyFoC39rVQuUA3ErpWgmG1HpoOC4
DMt3s/EEV2R8shorxgK5gUl5zjGcSpq5VtSWJmyi30zdIVPeFNVAS1e3Cvqn0zK9taVq/WHOQ5SO
WcgpvvV/lVxE3cCbeBUrATHzsPIfn7yrd0W+Cw+cG/02S2w6/GKo7g/HN8mrPv7CgqnbFKAZFtmy
pg3iuEEc3YWfRRfGAeuzmSYt014Z7UH7wzH4lAqy9Z40snee96pG20sIBu4hfchWt7UFNqp+kRaZ
VbrS+hCxbePGWpNjEiE22DsPzbRt+cZK6do6ZJfFKShkkTM87fy2MAgJ5+IlRsXKF+LQpqJSifFn
gw1PB+2RwlWq0NFvV5EmxHlxJ6RH8+exAvs+htjYv1OTlMV4CH1PA4sk/sC8QBy4InmAb/o+x6AQ
X0M0IqPAlWysxjm5fgd45Fb+ID/SLtWpBRXfeBP9h5oa1oASboDXZcqpwp0Bu6OHeWFs+wvCZOtW
FEo+xPOXLL3zPcUCczw0nOZow9lau8fdwKwvH4x+RuOyJovtLhL7akAWehyZ0jENu0AYCl1FJDzG
rSKeoGTf84CfoaDtwiYrFi1uZW2AbETocNbZcwaAuAvJyVrEqbRefoX4nzguF6M3obi8ubVhaGo0
AmDcnGPGN80YgTOtOGvIKXEuFLJV1JyCnqnJO1vFDejVa1SU2dCfUg8/WdkwhVzyCxuQ/b3tecKs
UGLweKadeJXwRVwk4mklu8yZ4GHVWZXX9SvvTHzcB86UI494GleVDUK4tYhYc2oMFmgkaJJUzQZF
ch4bk1cTVQEeVIRI0FbiyI7BduAKLsJR7Fcv48ybZ/XkIue9Ilh22P5lj/nhY5DfVvYRkiaEbylw
rKkyqjLZ2lm8KhSPq43n04dNOyWmJ8EVYaaRpv8fWf+g4goNYVtt2UDo8QTWZbDDJTQxD+flhGNx
WOBO11rCvkGHl0q/YLD7u+TGQaWKUIIEVJlVgh7aqMYoaCnPe8KtGIMpomqIwZdz8MoudVO/qaR+
cnxZA0kTBS8CfNuYYITXVAIENXwxKOWOcfoAgDvHdQB32Qk0kBa0NDErjCAo/jvruRizemOSUUtY
8pusMkCI6Dk33fDTrtMvW2Nq0eBivnpJLbCekc0nSVl+a9spSqVl8ZC/EnmL6aJpzenm1AKd9kB7
SJKn2HthmceSH3uLXsa0KXRttHV0JDFxgS6toLSWw4pH+8Aabz503vna0nS282mvg3ZyuEEjzpvZ
hPI4HHIBOtEZDp/nD1PsQgVdSzL436U4qOU4yQp+Jzb1VSDysUJaxqMlG0rF/iO3WMujgaXGgb9w
0ej4oopOmxHk7tsCdsM4B8k+UGkobAi4cAkgPpxf4eCxAQ7313Fv9ZZCDu8deWcw1+ALxDuxwK1N
1zpJNwaPJddmGlV6jOXfsVYXunp2dMSQmwm4J5fJC6D6SRaJJ+el+22C2O+J3XJjJ8C6+DO/6tng
1oNu5M9C09PgEzATWuES/m65FoPBXHJJ+Dkria9k3xKWgp3jjadEAPNwhx1MlG9FPl3rTYZdWUUh
Ef7V49YH4LnFoRwOFANPcEjBiMT4CjClIZcnHupDAQhKir7HJ1YH2ERjR4UzO8cFz7xn3zQeJeAh
JU1NxwvLusfhsT+1ZBKEg41yQqoCOxBTLXIuKNB0BI2GOKOBNIMG8cKoBCVP4EVqx7fjb0/53LFM
i2/3g2NCqix45suHG1p4Q8a09OwCPSCJEANex7k1lV6KRePkp/KfKz0nR6Ck+7FOSWvk4rvQPuNW
BQcujuUPZIzjqA9qmeOTguo7o3jHzIju4TpP4KYBgkPgSvuHQMB8Qpas5xldC+646NDHWOal+pst
ETUa1nqWXCjL+OBbQg+dSgKvULH85BOrtWOtZAlj3mo6TNwEgeaPrJhWMhXMBVdfvKqTMCVy46m3
XGaUcjrSFvwMvAelDUEuUc7f4wJW0vZQwLU/8V2Lhb5WPhbCpR6W7kpHtDIqAOgv1MtsNR2qArTM
tkZ1bThTjf6B4uNdtD1iovfwxUp7eJa3piuvaPiJTLonjXhS4ZAG5Y0/GgJcOHZPQOsUqdFr4jVJ
G5h/p5qjAogzclfLZK2Va2wc0OCsVKXnNs69v4NJ6fCW3QzM5ShUmEPkuplZG0o37wVmGm1vvU4Q
Vu2JgOcNgAczNnc8d40iLS0qEL6W3cO1z11Cn0GN7x+zp49Is1b/V4per/3C/8Dq3HYmUIG3duXp
A47KaQiOXMwYlk0tAuNo0LjAESJNL0IFf0Q07Kbz8z4o7pmM6fl56yl9QGSOLyJ8p0aMC7Qs8jHr
tXdF/C40liigbV2Rlsh1olp/BsE0MVhqVBNfsY262diOoz+x6InXZ7KavA7/cEWZx9yA2sm0lyPB
1kDdC19pEbQcnIOWiuyWg+GMz+Cm76jekcJPhyyL1n67HyNRU2iSsKO8Eug2rQ9WdS3XBQa8BoQp
E1U4BGYYa6ONO+WCAVg2MPMUk2r6vdMyF10NoPVlEJqBBeE/21TImrgo0kset5tvr0Ba0yqLejpX
VzIXNJ58jvaVkQu7sVP0mcwtH8sLPfr8noXGnGPPbhJgXpG5/zVd7xSwGQuF/xzLija0B7HbulHI
2R90mje5R2vqHnytH2ZY+P+QhTN6dQv2qKpAb7+EuR07WACErb00NFm2xjdWf3qQSJL7IdL9FKX5
jBDT81rMblBnikKDW+Z2OUl3++3jKSbgKIwHzbC7lhb2+9NYg6z/GEAb/bHkSnGyhUnPI/ze+FAW
OyLZdmD/eJhm+8D36qBcBDmUuey2UkelMiBI1xY2L/Cf7B1t8lM5b0KI41xvFBkL50zs00jUlIw4
qCFAMFl6+lT7LYb30/iQ45tKs0wXijplYpufbzvSNWJ5+fUXfSbSUGNFHbQAlIzRWlfPY914+w6A
sfczkrEcQGrXSINNs4nJRiLf4MHOR1y9GrOGiy8pQiOl6qqZOVOiyvydyfLLqg5mQzJ5J3r5uu6F
Ukwabia3g2zYKU56nwmZ3uFdPMF98vh10+PW7JoOht3ooIyb5Ruac+X9Giq7SYBLC+DYV5sPiZak
3rNPLHM5nDvxM47BboM6KglNCDGWndPyxh21IICZXDMeHQJ13DEsyeDkGfSouqAu8Xx5oA+Pw4o6
dzZju9zlTnY0QEhimUkEjiEOaYRW2zeoAf4jNBnc0h1hDHSHOTuzeOKfyVoT/4HHK12cHsAoiUU0
5tu2jYLxFcWmj8ACLmHPIaQWOGzRUZQDIrhybUEgeJ/F3v3ohE+kGH7vJjz0NwHy0RGmghx5k7M0
PBGr9QjxoB7g4Js0pe2zQq8ksWw0eViHmXTo7vHnmHOAYGbUfO3IkYF6hwNigR256K+J/gJzgGPD
+ZzBsJxqE28pwtNW810evuqXeqEVrVayIw/kZvuH15vjatInsw7obz3haZAHJ43N6xA84s95M8x5
o6y3jz+oES3udFMAalqwxylCMCysKoO479YOT5EhiuyL7/kLLbI2UFHyR+qPWi/OBBjlDaS5IQl1
nXjWQzWW4BKXyZP3QKVFZFQZf6OxwHWlEtjDLVCQuY5PsqgSx44FPMNzZkEtpn//RJAsGHpVu6px
T5GQ5PAG1+LGqvOjQ8RRX7x4R317D4Wf/YY1X+gBQqmthluahStbmzL7+WB/Vp2yXE6LERvieUAQ
EY9H1X/o8prIi8JejFTD/977F3AwkGkZcw2aOTjXptqaj9PlbkRQICNMnXrSedLajyie6eDARaah
KKhNB9U1E+ZLSaodR6zt3GwnBGQ8TxgpvDzT6vm7A9Zetjesxu+m58BwKOdRUbc4JC2qrP8S5MxA
C9wsxJmVpHx52HT6id+7N7z9Xu7aDmnp6MLkRxIAFy4HrZvwaUamp1PXAZP+I1M5zpOt7DuZd8uK
FoUBl8NZ/9CyglFoUeTk7m9VPu96Qq2BYc/yCRMOvLp1752O36EvB8gyfk9BVzghljl4yv3P87Dh
8o1bee1DQZs55VbsFTiP2t/x3hszI55/NPBdOzEHcpzlR2nYM4ilkqsUUWwm3w6qAwVbPpC70Gt8
LPlJIiqcNownwdQDBnBoA4BJ09DgHlzm9Kx1MUypWldQoHh5fl9l9DJr374LxR7vIo5rCerxAgDx
4CaCU8RlIjuNfP65c2lZFWBh4miM4J9/TRRuFzhzp90v+nPPTusWOFs3pojUitqbeKrOpR0aOxFl
HKOBzs4Sfx93bgP+Ck2UX8Bv0EOIVTSs5afOBWtX4+V/WMFB0t7fTQLC0EqzSJINFlV8vv10WPK6
Rkl5RjQIhZdua91yMmW/h3ErGCnxcofbUp6p98tRPMukWm/pW6ELbi6596i/qB0x9ZlXkuVhT0K5
ugdL7DxrCkqzlGjoG/SP6nxN/l6kZ2P/YVEkznEhTJliIkoll9MVXE3Q9JXdLUhoEaWDvJRiGouO
+fwBBRikJUg3YWqs9mF8U6K0ODFpWJ5K+OEnyO6UNbCCr7uIuh58vAx9aRo4pHUxq3f8iVFiHm6M
pOIMsG4av1DZQV46UcFDGFjJjZwQKaIHHjD9nfBslgALHzCvKlZUbkJiVPjP6Jz8IS/4SIjwYOYQ
erO+rFvPHuj/P5UZ8dpICJFgFthUx9K4XwFZ0X4wyRweLV0Bauxofii3Oy5GuKuuDzskMVfgRCps
/F5s+uFjyMl18MgveIF4ZCoWl8ffXw3PL8D+Wokey48QPQA1qdyj7bgjZn4gaOd7lMO33RlUPOAI
wTUMsstLWH9DJaDMFXLI5BWAzKoKvOO2c4nzmEHxasMLlqfKdTt65xDAGsRvw8IqOUxwfjSptiBg
p9cpPBKTkEFFKh8UHlxKESrf4pC5JKhluGUKGFXFKcMWJscwwbDLU2lgpsg5VGfd7M59wSg5rmme
qgrE04h4vXizGAkSmaKI7QQ4DgHtNIh+r6tB5qtm1BCujhSHV8kworVpLIeq+Fjm4+MBV5bJzTTm
uwegP7EEnJxALDfPnxVM7l4OF5SFQ2UKCl7w723VAbmwuWYzBxWSM4qmqQSXTyrtye2iH+mnO8a4
zBfg1vbiyvcchK7WSoZBflt1ObFv6xKaj2dfghw1yuMMbdRr8ZlkgKoHaJVg1dUJfTnjChTWCIrT
bUCsG4wYfbu0PQmW3OynjSGobnpUWmlkm630iDWp/M0uZHmXPX4cuWOYnjhVStUokktSEiNWSk/+
Wxdk3jSvX1iGZLihRJnve0bZRIISFFfLYFYfFPpelINKrFVOObCpgGZ/piu9p6Sgy2i6txDnVua9
je7blXSdNqwv5u8x0lDpDp56vrNbwGlLxPy4YoBEwZJlej8JpB1vHOwfV1Fy9bUu0JI6mw289c0a
/Sc2GjUkfeXRgIxsrmj8r6PJrhdug/k815qKH5qgm4XDrrLvFRHdJ/sSejdJIEaSv+aplkphzvoE
2+fAJSF6SjizhtxFI8MML7vu1O0LUsvRB+xf2SQ7sphk4WL3ccxCvPt88n7PmTFrSL0ZwF72IfFa
tsDCukBUteavBj/KrK2QIFbxrAWe7CINQ8GDMLsTFmN/O3EdT8YsIx3ZAv01cBxRQmltbJav+OLd
i6HTo9ZADWNOlglUEdTG9y6/J7XLEL/l2Ow0xbAACrj5undxgmYheADzru5dpjKFXfj1ppjxFO5e
v5Vq6Nc/2o8D8cdHIq+7eU2PB/Y+VHQwlJv+Jbgfuh6v1ItqaEfQp1YjNECEH+WsgQNgJVDSU/Jo
eQdaSsuK7UzHmou6Poz5xgXNTRHnzMz6dJTy9EYtP3VxwA2vj2B80wgs5INP83qbh+RlAvsWkUB6
RWExkb88RAh8+f/Lo+TsA3hLVJ4LbopRloqtQN+1g5OANJQmxVgO+9LCmQ5jwkNcTYGRBcuxrEm2
IcvI+L4jTTOP1Yl7YuJyruxnus+s2aA+kkMltS8vP1Q2m51nwHQBwRMmV7OCfWYJv1ONCcZt7Fti
nagsIQ73VccRli6m2FGfwIgDpVmi1d5g8CNjSSVsof7pxcGaPD9u2wzAnpyMcoUUPYyeH/tt/voH
r7MCRgAvoeKx0XeVGkmVS7AcKNjZZRWbFBTekc0rWSr0sccFI6lgXMXUU6tGrg53A9s//lJeBecp
YqJ4GykzrCFwDxdWS/7Eg/U/rD55zFirDsvTvekYZ54UaWkPej4Ce1Bj27Rgqhv1rOn6CzEGX3Du
uSeY57IhwrPeYdTteZCexUxztNw8ftmo5KP4EjvmiPG0rfKN6XVRRVQdgzqqtvzFaTQR3q7NH9At
9xBofwZ/gsoRdhQhZ5S7xlnI6UtoUUfc4QZZDY4HVnBmMGgnoKa1xQpKlahqfGsdJMLStqnyjCJU
C9rs74RQND7bxWepiSzu2kBZGac9cGw9KSV7lgjX7PJqa7kXmPZU/Y/RY/l/k6dkF+TIo2rluz9O
HxM0hu5V+kcJGdSbqGbilWucLJFuVxhf2I8H1SsFHzZ2wHJQBQGjYC7D13jPXlAJAHS7tlIqntHD
KtYR4Xxlwa9MaRf/YawHhwDOgegydZmnamdsVd/tvQcz1hCckAUbbNP2ZGWo/FNtnWDpeFKZnQDe
gtdLWwHJGSXCC117NB6/jbV6pvPDfk2tlFuIzbODnhaU4z6NV1LOE2ZN7UeBIOpxtc/NLxK0H7mQ
oyFZrGCCYiHgY72SxgTbkGv5vWx7kKd69b6ps1EwSIOKR4bZ//Uaz6rtdNRRTHixKa45Tt4VzkNL
Xh52fN8IGMSxPc6VEfAtSpe5J4UF/9j2UVCmiH6koFufkppKc/gFmikb4hvk/+80HrN/GlErc7GE
FotAO6DvXslN8a81H7KuQk6MuNLKbwB8fhpjSBQ78hIA2dmPD9nq/TxRokfmSiXPsrje7vGaQFb+
14KAkPt/Pzp1+IB+vZ+hSjtadjTKDwOz2Ua+vO5z9zXDM6eNjROacIOfthW65BiKMoVID7GNcaBZ
jBfJRmRETJNbnyzZ5vynsF+DGb85u0eGyfwHP+NEeU+5P74MwH8VTGOokatYd7WgqYKBXnDcfL1Z
CIE9QWm7fBP6slZtwUFs14Yr7+sxO/noQuMwBGqM+QmMvBpLjFHp856/c+YSqzam5lKZvidRVk56
Cy62twRdbsxafpThUtz1QP7gBKKZtn0Jq9C5SdH9sQfsfjYBT/een6dd3Cw2bSKYz1aP66VNLE2g
YNxVBzdJG4KEBiW2zb4LYkdPMr5KQLLfFYvCVM9fDxiTClFeIomvzwMWI/VuCtbvuqkiP7Juev3S
Gotmy3d94t/edrljSddiuaxMco+/dWK+pSQXi+h5N7RfRxLVQ8BYBYz/5GKBfLYeFW9b7/zD278I
IRx4xcZv2eHuNztG9aePiLNrFIavgvHJbGSsLhPEyqEKZEVy+4U/xKihfELP303xdMfJmuYQhfjG
ZJCwttAGCOIByti5w3LHcHToe0W2uBCBkkGl7AVpHOrgELNOWAJxzCC9tfPxM0M+MniXZc9XCezu
EH2S6cyDS7bVzJXK5Z9v/bOfzXRF3UY6AcimYCpeaSWat7T/RCZ8+i/wq7pZSjN/xVkU8kiGW4bA
jrsoHPfd+cboPnd0y4U3Q5tvip6VFx18IkyJSfoVSBxBYlUNyiNkvt4iYjExhasHGHxhfWDMBmPY
Bec5DNJEUGRwDeE6NibmexAaIxD/jA4SsS2TQfPwxMbUX46GL9QhToQnLORUizEDsDLPKnTd+zv3
pT8s9wfGQoWmQU51bs/ld+8pg/PD6J8dSe2kj4PG07rdi3kD1pzB0iiH217Tc9G//sLpCpfF2NZt
na0r4q2QyTLtlz3jx3wgiG5D22Um1pPD1h51gh9RaAoaR4GFKDb+61iFENK1adizs3RWx1YDLq6W
F3DMNYGADW7dIlP06RFtpvELaX0r4mr1g70quAAHPgAIEj2MCut/6GK1ri4+lfbHIVm2RiSLWTO3
scjT6PAvVdLIOyWDSzpvpY5MyClpAmKfBCd1FLnHxy9yKvvSOClBtqJr6Q1yXgDyxM6uUxWS5GXP
H9difhsUgkcmqzB6kZV3BBOrRNoHVZ6XLkOCCVkwVd8yyI5j17TErRyCY4+LqgdJ5Ij9QvREXBvg
YS70l9mEL85P3EQSuBlLqxDy2Az01x+Jvusy1yuKrR5fRRWHTPT8wTqCZ3pK3Pve2mPG53pwUs5S
/1yJkN9FM34r2/JAFG4iLoljsFlB2Yyu2Ruq4HlKG12XUEijtYES+PyUdWsz6E2q63sBzOU6Llnx
tkRaH6RpG24W6rDdyQJyYVutI4oxjG4o7/L2Sf8WwaQR0VAJF1Cr+aPYlwcu8lqGg+eosyNT7LmG
MyBX/1pu37bEf5lsr+Q9+DcbaslSzbDlUuYjLktv9cQF0EPRU5SoksJzWUjyCxcaR7YvV/X+TSpC
Y2sH8vu14wZdGFCnlGAFZGecek2lE305f2lxNZKoE2fT7Eieh1M+bVcBBuakN2z8FhayzxvkE8wA
15CJCO9pvi/Pr/hTF2JFbV/lo8TBSvr6Xp53ztTUNWGcoZJTyGh46BcP1UjLX1gA5o36inr2EIZu
AG5pVs4ypoFC48peiOrGMTAkw3+0R6PDSvz3rCogdUI3gMjZgJZfHY8I195ol4IdaEz2m8mE4vuK
8AgUjDGKp4c2XM0JC8y7URfDuUH2zyqtXCuAIPCDHDO2zFRJQtNLl8BJDny7MbfFK6w7t/nP9Lts
vrrakpXGyEMR0ZJi+7nuHpDq/weouE46xA9TVyJLpfxjfCrkkwYZdiHxZTIjHD0UV3fYtA5BmcnE
H+UibKYwi98xZHbN7SUgzawybCnDb1IOjxalZk39qEOW5X6b+9adZ/Y1H4Ye4hRsYZ9QRBn0qAqc
8OGI14xXE6OgppYGlVlLE+AgiFCTsEjm/8Jzue7Ymg/AdKcfW9fX1MyJcHV9oBiggL/BYHJaL6x6
c4RaTm57kMt/0CC/d8IdEC12DnZJxt0o6q0VxHiop33NAiRQG+ZVjusgLaHRA3SdAsXz4C/XmByS
hk9m/bxHoXPqhvDNag8KZsVnV5bUPSKLqEn7NPmLwEe+gRYVavI2m/AJ4X1MzEb780hTdKdsKSNN
a80gIOc60tLj0FNagNSsJLxQ8ZPAmwpyaSlbaGWNFSqvpmWJmVyzTLzmUwW+milPxTlQ2XNlTFkJ
Byt/eaamy1sVIdbyLKCKp7LFWeb+jGENGkeEW8RUf/y2EQgCe9BFYu1UDEAbmr+4qA8/EDy0sOxw
7AIuZjOtiNOj3z632oBq33b/rfnBHBgWkY9JXbpkTtFWBNnmliAysWSGOixdboAnGcYb9cpyNZ/k
0Nd4JqzKq7ZKap/cD5VeWDM5tdgdjqkUapfPay/J4Dy11TpQMLae2vW9sYL62IpwsYJ8+56d46Ui
K9Re95H/0qBbJGmc95tXMK6Ze62Si/jxKk46htUWay+Y1umb7/g2E1cn+FwAcNSR44zX+cB0mNZ+
e16t4MdFFbdHCsgPFjNLck2JJgURKOui8xfl9KC1rF4MYcERCIMd0iSIsdSC2jOStf0IxvzU0Awg
o/jauQxEoLFDLlKbbVArovXraLlFYY2majBBGpvIVf/mNBdiC32KngmXS41I6BaMZMPTtWLEhwCC
/gxZzcQFgdfRJJ7fJGpt04BJRCQ1DzVb2w8JhPqe7o/g0W57Ct2SeEI3/7qJmhSLfo7KmqQ/Zkm8
jUcXnXOia2gT86EPTPWPinp8Gljdv+uOzlpn8mV8ZfcUr2it0QILfhSVb/ITNRUgNPU4LCl+V/IP
liGnzGnmiqmDdGq9IfXmKunnUmrC7j7yMn5yonRakqAttQHBg0QxH3/znxF+Ejg07UkoYe6AvVwN
CHOuxjqAQCxtUvWoyXt0kM3R+qUzhmILQnRgTPvfLcsmvE+RCM8zdeXfFgrf966JuBl58xjQymd6
5Yyp59rwGj3ttpNRcqRrH/WlgLgJZSQolN1ar5b9wfbIXv9iG8GLv0jJ876hDbOSF3Wm8ZIbYLdm
CWgoyw4LHHeZKBzNSf9COxIhMdyHXJi+i7FOLd0XIkjDWwJCE0XEd0nghSr5PbnZPNk3naySr5fa
3tV+G1acdbnjdK0PR4xxyM49xgjNw4T8Fw2wbjtULztIyzlKjuUPtU9Tt0apktosTJ2x4uZ0R4w/
/I5WNdlsZlh/1YXPer6D12FFqiIrvtKLQW1z1MQAkHp9HN3Gdu+nhIEfAtgR5KDKA6xHvDj5yrxj
R3pM6aiHFgewLg2J8E3OjaDKR9H+Iw4fjJ0jWzj/OerIiaLuYlQGhgH82laJiRUQ6Q2r/h9kQev2
ZnrcpJw/zM/YwRlFfyWh17FZrcmbAkM+THxzdHFhrhWl304tdj9scZvZotLXc8vsav3oytHf/Xga
WZ76Ggo+mN1O4ANhD3qhoYE7tAPQITGp2Knk6qoG3XspdYtTajq9sLsk0NC15YAWEIGARRaT6EC/
RX4iYFd3KLj67N51gK28gG7SjRHX28l/DCgVVO7srGtWYLx7jSOjOBG8sBtr+qUT4yeRanCIAEnG
CqEDyujyXRKyVq4UgylfZi8SsUnls5iwck9b6a0tCnCpLKkCIG6qEtY3xFwvX7xcnklTY8YPyWZ1
0siZj8wnxJSK3yfbvswY7o+Smm43DWlwVw290prnFf0aEKpujNvxoXFMyXogPiSAbXb/Lf5k9ndQ
Ok8GH2DDPIPWaAn5xHqV4JM49f09nxQBpBRirIjC6hGh2ZVx7hFTXvhTqRi64k+pHpgQLaMQ3fQE
TvJWmy0i1487VyK01/6V5yQOYTbYa+BeSKYW5Ny2eTgRQAwyBhAxqG78SoNWJTnBGT+tfGYGtXOU
df9JPQ9LsaWnXQmoOcXtdrcKLF0A71qumSx7LtSPzTGj2JUR3Q2x6QCnq0H4TKzCq579u4t1J8gv
V07CBzHLraDZT1c7hCTDFeJZrDU2mHTd6mBBjhPqiFDRHIZtv0NPJ0RKrnT+PCFb2jzYTNYw/v2y
ISSgLQUZ93D+2wxKENrM3baOmeoDEtEeyy7ghZrTU5ZdVUDrMriZwJxujAb82AijNnwSDor3LN0P
wcaVV3LPk7qqB0OL7/bmBDZllVm+SNJllYj2rf4EV9vS5MwjSa59nABQ5Hofatd3zZkKKQVZMY60
Prlm2qdenbGX7DrbtXGw0T8+VYB2bqMPobczIf6zmkG6IuIxBhJL7VY719UqjOlp1gFCPNqxv1F3
/okjjA+xsE87tqUsGS592W1wG7aiEFjGilYjJXeol6XJPCKvEiwYGbTFQ+lIVDZ7rDdGulZwjoHj
VIa/cIPxYEPTYXzTUH5+SPfKKO6fS/4a0vFnZprgOPZwfsvbhRCYBFdU6/wcxxTQfQnyJuDV6LNH
17sPrNIme8jwaSyW3qahO9CE945LIEFJwwZmVKXYfEVCko5uB1R14ORZuB3ic7nggUI3UhdzeUyW
tnS09ZFpxJIr5UEOFh7P2LQVEN47aiCiufm/OBHc7jLXT7HXrdATWKSX37YLbuB3iXk43qpNlDzE
YaDRJKv4t3gO+yQ5MdkZgYMtlkaPvkGyU7cH+e+40976yFyfzV3e5sqyLDKU7P8MgpoMIOFx4bGH
8nDTmYw5qG+2OPMrTWw+hQ08TFXsw4IAuyeOE4lu2J8ljBqaL6iTlKcQr8MD9SlrJZabyM2QBvvv
46vyRBfxmATv1p150cXGJ7hW5HjtJXj2JNusjr/esnrMavKDXSjiUWzJ6x3GaptEdAMwivN0+YYB
HttT3j0+cWZJJfbnnxQBAcx2GYH5WoojRiI+9doNPlk6QgEjh5BHkUzLuF4rHEktB9z6Io06Mf2J
92tNvxC1gCpS+eo+/acr3bS4l/LdYLdNJKG5Eg8+9tmzFZ0rQOPGZq41/M0NO7QN4TV4+ypGozF+
nEbCm2JgAm7aLKjhPuMKH9uCTGtR6V/4/uTZgfC8IgE258GWiCSKl1N7tCCca1IBZdT4jJCjX+nL
JSVhRswHf50bBUuzUrwkDM6IlLVuBWknRfMJ28wVal+Qq5H1hMMpHYY4VTvfQxrJ6Q02k6wsA/Ty
pYasMmeo3OQCIvYMAaN2d3Z7GA74HseWxBw02GQ1WZNIVrZ4pYtZzuBiypaxdLwawbpdeH91i7jq
+rK0MhioraflqkKWBrBxXuXK8BwaNwHXWYt4vCtSjjuXnAxUWtCf26EEERT5pKraZvyXfsg2UWIC
DnRy8FZtVpb3XJ3jhQC1y3aKBP3pVpV3ApHPe2ufnucq/7ZqMBOCbgpAvgpyieP/V+PlstlXj9Pt
gT/ZpjquHl3H5TGdDnDJdO8Zcz5CpGjoFjBXO1SbgyOYFZUiGEIo5x5SAJyMaRNx0oCaxjnfuMj3
jlS5AHv+EgO5zR3lqAI9HRtZHXZrMadtgHxcji/f+FWoDWVnXU0pHbv9DFrI2Xk8P7DyTJCIbFK2
muIJPZxQwLenv4BFNyjH5y36jyskwqmGq7bhccqNzjKq60qyiCWo0Nj4l328L2IY0tfEM1vcEF8W
uYwpgxrHMcYn3K9t+4YFxmTy6XxNdAB/CP4uwckjKYcW79iCeHazxLRmCBcFBf4S3WoNqdB3s2we
DAq8bzzAAcgSqTTXbtdLnzhl8lUmVXw53LX+w8ceqTENn4lu2yExL3FI2DTwMK6HATCVbSQr1nU4
OJsPZeNeJr9MeQ85aDsgyAEYxyEJOn6DQ35Ho4GmeZWmFV+G/opOaT0ylwJpzMM1el30jWXAGRBM
c3I4qaEnPIILJreT2zh5glxCkMf5Ttx2tlCJ6+5RSbxnUNZGL7VxsQ8z3ZYpvYXa03CiU9nwi0cL
gJksq9mxPWXz37D+XTrg5yu7Sw4pJboqF6Of3udkXN+zM5iBrk3/vWWySXrKbt6wOXmSZvseKIyT
ee6ziyfflGvJHzfqeU/NjTmW6q3quuPHRMae8fTfgeTM9zo+zdmpOSpCuBPkss/KN34IYKNU2FmQ
NCEQC+kSJrph8ijVouxhwcYyDodwhUpFV7qyJyDDEEGqBYyvGhqv3pwheXa6p9h8/rsHYjzWrBaO
Gmky9LlDLtqioGa9isBrNzykUpUoPyrjw1rLlGKoz08TzOyvhNnlpCMkCUOdK3x2uGA+O+Cgy8L5
Bf8sx/O3SVtjjxQT/I+gtbf68BS5Qu3KDEOR6WINs/tsWEboNrfJLuqIY5DKLulk27JP0u1EO7fH
tIYPg7LfTIN1uyFcL9OaKAkKTb7awUXBixxPhoN0jibc1Wz66pW66Oc652dHEgsPFpbUZ3DksUcW
RW6UC4qIMxQ1JtO06b/qhDnWGIKM3Xv9/ZtK/nniW+D/kOg/axWJJM9x9FHds0Lx8o1tzpR+bxk+
dop3HZIDft+QFlEi16qYebX/E6Li21+lV3YjGEWmBJdMxUSX/FqF53x0VZ7Bt0UxSxkGqofnehey
5HiGVVgKBGgGfD4TFkuqy3z91jnSIpmtNEpTHLezP5uZnp0kz58dtb0MAOqPAd3QYWN9P2lP0aB0
ReMiV1XVEMXT9FNm0s1LQtpq7FU3GyH2eco6mw0jTxDB8F13gOFR09YwMis66cK/wGfU90LegYGs
TTGVPZxgBJXL2+7xPg8USMN0E5ldXzTjjHa5FaZLHGkh8Dp3k6PX3r6Mh77XW2tAYqoaSdVBFfpe
Ko1lTwnS4VC5QF0RjL/riSCrhkLGimBbV1tygRpiliOau+zSzNepoSixxWUFabersHAXuUhwgIEr
Sw/zryLbCyrVdHvzFIktkeMsxsxQRKD8e/QPiVb5BIhbNNzUlD8zEiJhA4uhn1D+OYTxxvXN2KTR
UIYazYykE/e4ukSWRcIB8zlsJ5uwcb23zB/KS1B3o1wsKp2WWkpEwmBTn1HKpwQhnZPdQBfVJxft
gyFC42CVsoILiQJOzx/unmLgn4RUiWaZkb6BuLHtYHCmZlgFB5CK/DtZrgZSzz4faUN7PVIncjMO
hvfc0hI0XyCEzu8xjMLZZ4ObpyXNB5eOLRiTFGFbiqFtGVqob3CjUoJ3paMKqLk6M0fK8DlcsMcF
uiuW9DLEZZkE8Enn0RdvTy53EVVbQrEkNynuUY7t+lgtcMZu7ARaxSOS1xcOwOqhM2xjpoZN940P
Y67V7JHPnzrFuuN+YvRYRcEKJkGSGtJiWiRUV83VvIX4jcYdFZ49s+bwX3wYCalXJ66K9hA0u0gm
SJrocX2S8yztfNJuvTqCa9MHCSvUUTPDR1GY7jAJZSuseIZpI5ptkx6iL55Dt6E83uXbSotPVR4Z
qp6OAdEczp1vPe+p66RREo6+jn2Osh2RYGnt2JCfiovCFOKKzy0gU8z2AeeBNrRyFltb2ql/RJ1C
FDCpmglBPXfEJCp0p2c7YlGx+d98T8uRoKrsnkUGbiHXXfW/XT7HLAaSmZH5UuCziDPDWh7IyX+r
X6R8J8uaPRhj97lmxahHTD4Li0adfa6lulEtEhIRWHW6NQVNyWh7g6DFcOfhb6AtSiJtfmcWMNs9
Sotmsy/pNaftCf2sbykVOry8JVBjUw8UtHOqCYUeYZtPLi6OlXvxT/MlFEF/5SGPXziYWNdIO0KM
h7Xh/qcAbZvb/lBPEEAKIBUJV/HOuqoby0xYxLSFz2yL1tuuFuLhs1OBcZfaBwPP81djDRhxXgca
T0YYexX2PwWWL1743iUzn/HttJTyrbPkWxrdSX4tRl5HLbZzXpICWoCfiyMoZWZ7kk04f9q++3Ds
2OHBOwsJKczSdxAE6I+OjjCgAAAQPo4G659RBFUWQbwvxtEgHoUykChwUpTSyEKUG43yvG1SWNsu
nKDHeimMU48iGqNHenLoBIYKvc31xAsvHrS9uIMOVq/d7sMBYr/P1KzL0jJ5hFipfOu8i4lbMA/a
e3Syn/scGmq/L3Adub3AWrWhNV7QSxzkSgGTtKH4C4uoQS/aVOuXGNOJDwBdpewH5w8kGecC/Dne
/F6uiLll56+FUiDXy/hAXBAZrfZ30kcFQZAmwcI9h4BPXo1q6Aj8A7cdRm2XrC2PfkXl0TDXeYFm
gUvSa/+egkJzSy3n5IikrD+SIqQ1jK9/8S87B3VBjcDYdJI4Sxhp5ga2U6J6FcHptDk3W8/D9BHb
rArvl2Yb0Ot06HF63J3rWVR7Hn2iZYgFp9dtZ8+BfHzBaCWVaXxW6W0zIQ2jC9vvIAX/QmI9sfvm
MjMJlC78q6OIponG3yCsJ7DoQbr3uLo4bO9Sb4x7wM2U5PxhXYDbcJl517fSDOH9Y6/0y2ijid2C
PRDny1/cWR73lw5ar5dW9anE51cOw2oUVGbTDM8EqUfZH+KPIg5cKIHKwSs+qUBT63XvxiBkp8D7
ZI7xNlEURdMCGU4v/xjN9XmAMONGEl1hccZMlxxrBwRUClUQBF+iEqFY0WK4avV7XmytEwQVzGY/
Nbp4l3HGZzFNGfUNnSjVZQNC9Hi920daPDLBLvzUQW2n0m3TfuRLd3P60pv9d5GbxPKYHdXQrYJY
ymP39ZO3dNcr5IkAlst9hQ/nOOQgNOoacgZnrFq1DsxJU5b9ZCUvcRBGZ3W03U5obvPsriVcZL7u
3+cocZgFPs/pIlI4OW4ElNx1hxbvr2CbQRBhPFcxOd5ZHU53lsywvo9urTrQzbSOQdKxXWrwlmVh
QSW1+GRnxwYQ88DQ4Kxrq5rSzlkVYcod5ESMrRG8b/OoO7TJNiUsoLU15mdO1/Ux6KrpDuU6UM3h
lLHS1zZBBZbnVcc85IUDIzDfssBsyfDm6Wr8tHQjW/GdmhTI98RgL9VfwiIqXnyfRgZJroGzHjP0
BHoRGaDAQuazTb0cDCB7x84AvVRUS13axBJqYRSB/smiNzCcJat5Ta8mWr8vCI07IaJWaSb6JRua
it1fXtrPX33uozOzbH7G7Pq/hVpZjN5RjfUiuVR82j/F1yZosfgHKQ4d3sKhivkuJOgWX1Olnmsp
A1bgLP9yrHqIANvAYAiQGGOhgmb6CCKY1+w2nntOaJt/hvB8E8JganXnusMKf++GBCovm3hRMucW
2x+UiRAJsIinMnz//TlcZ1I+Op9AL8BYKu9NGg4KDlOQvV4yUL7z9Ve/IW8S9T6lgRrnLPx3YJUr
yW22GDtIEfrT/JiI9Sp/4xEZ/F0Xrl/bj/60xYu7b5P/3Yop+kDrmKdXP+r0RJzOnwnQu6bxUCjb
UX1SzqP8J6J6iIxslcsSoN3vI2HTuSeKvfhRYeCdBrA2Jva4PjxSfgzTcDVk1eUNOzO9fN/rnECo
jKE19yaEzH2URj3pUlTcbOzWZ+aZGlbrUoE9JEfpH4Qhh2SPzrjhfCssVlp9FRLjdX/iXoh7xg5d
3kIm3n6NvKWyGy+2UlvJDCP52IzbXH6HXHKOsA72z09Ka/LgFGixUlzuxjeddJ0txT5HhhtTG9NU
OWTCB9cHWpPDLXkR71z11P8vQv/bunIipr7lagg/TMbYtrUAHbCtLeS9ikGMc6gDgk6gwStBLpcS
0RcbYCxRMGcRnfSvLCs1ZFnoa6GOBogX+0j5/6WMQ4NN5qvvNPEpb93r52uOOlmtBfLrOsPmDpIK
86gSlp+hFzUMQmz2a/A1kZwN6YSxObXj7WeIVzM+oVwEX48Y7oM2X2VRYY/7u35DPmeyB2PlgQfl
pKGnYzxKs01G/otUDq1eHJuZLHw8V0c1puLXYyP1dWkGvm38XiRxdDHrp76aNfH7KVM0nSE6jP8r
avik3BNkdqocNuh9tJikngu0aJfM2eNM0KefgXBvVS3Nqx7F9bqqawSYEFeA3IhBPZpuSBhb320U
B9cizcfbwBr81u9YCbY2wzVqNDGaYxIikmFgFjl8XelF+/NkbylU3BvmVm+VJefxfL8X0bImWHUO
7diq7XpsBn/89A/7sxwKo5447hJdxxT892OtlOyZD8norrnGF9IB4hREcA8Wy2R3qQmDE3xy4SMV
dDq12d5bR6aL/d5Fy9mSd4kDb97kXUMuGW2eOUvr2M1j1Py1k4AqGqlaJs/oz5RXY3qImtmfw3rz
t6yvYY9dp5nucQ7nhn4gOrvIgnJZRMnkUgXLAhYZZQligUijdZPDFYvS9ZIRZW3jRYK3eY8baba1
hBaSKeaP8f04OeNRkubuYkl6ZiPMmEYVk3gNO6L84cNcMNf5snfer5aZKTSx7KSCYPx7XHUrvhKd
bwt03b4Gqz4fFtl2s+ew6qM00JNDq9JxPYprkHFI9FNeRjVEmqBddeyMVQbdf8Q8wF2OOE5CwU38
7DFlM6zuDB8Gs5HsrxPFemLTIn5doVXZWymuevqj3313LatpdPZEo0ilWlzFeDhx5tZXRS3kbR/1
3mPP2EwVdqqzlvjdKcx4jev5zMFF02D9rnJoPsLZMZ4S8htNGDJYOShi6bsTUgKBmpI2JtqZ1xRG
5gkR4nO4lToO8MbAbLbwamxYO0xkkGiaeptIu4EsW1UP1EXEefCqYgMLVWIPEbUE3QQoidXPliJ7
O8XBzvtr+LGvcpSgIdEDYGrDEevCMGWxHFraR5pvWx25NVG3eu3NAa74gl+E1HsGU4UKGKJ/YnTU
t9+oxPH9Ub4KXUUgm9DdpWOPDQ2XFejfTpVg2SWLIPH9e1GPj9ijcTwoePLNH3Y2uxEEWKxQScKR
NownRxIKItIzbsH+FV871MEqnNhMmXxrQKtC4YHqhF10Te/0keul6mloTn4XP7TghcYljiK2zc98
ylxeWIgb6u+Cu7fDiKJPKqT0PJ16ECE0i2NHmQOZcqop6QUeXw/dDKPfXs3nb7/RufU99PxtRDmo
gm5Ja++oeun5JYOhr+ppdQZsu1tquySnRiINwG3mn5t0ib7iaJokgB8+nPyHSu8Lps9Kvd1y95FW
RSXS0eiQBe2aC6/5FV/qCunMv/bU6vkevZwYt3s56iicic3eos/zJrLOIkruNK+iYjbM3DmCWRm6
4nsEWhpbzBmzxGz9QPBJnbNsKNugZHC0g81S1Rsxuhjd7b2lmsNSpUsDu56qO7Yx84QsFw6+dQRv
YmYqtB0PAmH+q1ss6cKPFYtz5qhjN3v9+gAy4RS0M5WBqPbhtdDsvexl42fYBOpAGrI/NDCIhHAv
MxwwRqLonHFxCHPfRrCUmd/+iCik7E21TzHTpkuXxEkMZF2hqkI8fw/BzkbH+fjNq2OL3sWYrZ0l
YJs2FM0+gryg1j+mSLTNF3Zm8zIkG5OsFWF4k8A5RDN1GBjm5bAaQnSBjvQv1NNb3vsAqn2q5fCX
BFkoFOZuyHDWUjCfhPxBpLkbeGcM12jI496XsNoWffMUqFPk8GJNkF2d3iDTBYERPXpiqYcI8nMG
KaxnehjSqcLCPPR5E23GpD/FL3vhgkHOXunKfh/oa52EqhLwKS6Kn14dcX/Xd/YebNuC3DOyvejZ
Hdv6JDGyrPWFLHKe7aygIgcJiTxskvW0u36pwu4sjp+o6NmyewqwYp2Bnk/vSz0YdBw30T4Xb6mF
IjJEkN8g+gwn1nFtJOKZwZdk49K6LNwGph13mz5mJNhtwFw6mZ8bu19q2ZbswXUA1sAnHMrKbBYD
7ORtU0mQXLLhpbmDLZajZ1BgB7OYQvbaht0RmetnZuyalIdoU9cUxwhzEwA6P4W1nKR7Qb++D6RQ
HpP47qi5P7ymoggUR6wzTEWmLw4OaBCKgQTOjlIKEwiDxzizt6I1fjE3NLnOeMulZeMZnelzXVPQ
VVDpUDYxKjWs5475WAqCK2zkgEQ57inPT96yN6lfzqVxWhEXHlwPa4xqhc9x9SYqSoHBKTYnM4Kd
RfmTaKW4b+RH5S/HstoNBMtjKS/ROOkklxIp1TDmxR4lVS/GMjGcexynpfjJ0MiSQbuNkjE0xN9c
BWkV6+Hb5vwJo6GbELwdsbQmgRUJScd7captOoK3VP7YK9NnsKCpwDzIzSF7gcwSMiJM46Fo4bb4
bqLjzK7ZnLim2bx7UJTaPKojJVcn5Cjeefhx6KWSqxeA3lo+ba/685udwKO1c5H93BDzp0A0B/PV
rkjE8dcFF90occgze8utSQB841IJLnq86grLwJSYOrYgtNQVHOgyfPo21iV8pKVpbKDd/XLKPjU2
cwMo/dnrFfwu1PHZUsWt5W9NbGDy+U+zjCNSiTOJl6J2MH+Sm5mSwjpgUaxl/czH9ce43kxdfEPJ
NAJlRnR+jVICHtk8PRDlhaGt/Z7TjsKkQrymR45S44td/iaJF/r50QY00mQ+VKH9wwuF7QXnbrbt
jgi+B0uWRZzZTSTd03mvCHc6wM51ehixODro3F8+uOWYrXfMrHWl8Ay6J5IGhjdKUXIZb6LyQpI0
hrj9hwzc55DpNCopTvIjFofgDazp3E0Qko2lw9g/Cs3utzy0iwFTVxwyvE7p46C+jb3r/wfow9Eq
N4vFfgSfPuoX4wGH4Fw3PvSIdj+gRA6uilM8pjALYJ3LxIxE7X98KkU+BlV210SVAvC2n/FMGsPz
qDQm1Sf+q4BYe8jrv1Bkt5V8jZIVa7UReqj5WY76SwWjIvwLLe5rbunmDZrILWs128TABqdB66OB
gY2QHyDEnZ27ysCb0aXJewKE62rvC9ADDt/GKWFUXi3OERTNIptHfXmCoQ3QtBYViGha8Hxd9wjL
mX/j3TpxPwBRllDHGEKXwF81nGJ6wpQO+DIHFe+2cA+lCYaffms7pBjB8v3K1EZG/rvr2RiE25sN
Mrd2qPS2yk//SbIAymxkOu65DJ8wR1iZOTRVnkj00f4RkHa2CHjr3zZJ4eiPrZy0FDzl3uMPejLB
H6ofkEb0gMxwCgtUTAOppsAnra23kYBNCAvtfq3e0JTVEYJ370TFbRj8MCn2qiqWnt5c8uRrvff7
ZxyHSwDXWmctVqbhs54L0MReqjtrP9sx/BJj3yiyPjOHZWZ+73Lh975uDkL1kl5FpdoHFYMLgcU/
uJjMLlyqeyqRTlGAGd9rb0oCg/EPD56GTD+TD4o2KoLyjwnM9lcDC10fbRB6nYX3W+M58GWo7Cag
YhX8a3Td8bjrK88EXqrXuiOfC4iA8TBFsUV2o0mB9iCOU1ncIXhO7HkTgvruMSivsckQxb3jfhXM
23T15NZpjaQMJdUSpNrgWlW2F1M7AbdZh+d5TYtnEnST6ZC/Jug2jKx0C12pTGICtVzM5dcls7nh
tfj1yPiTTZxLF1SCSJ5VouzCPrhuV7GuL7OJBpgQLG110A6Q3sS6vYIhm+u/az0qcU4lv34NdOCa
G+lzRkNwjHUE896sQhxzVC+cvq2O5xuQnqWdOFUzeuev/hSGExDFlckfYCu/NLV7UG3dSw3Dc2wY
hyrtATL0MjpTB+sT+O2PSc17/dVfNPlW6ng0wi/5njZEdkUkjdLHvPUfCkwmMJoUDDmZ2CyPqa+0
7GXwTckMawRCc4uqV1/z9t9qopj4wzYwYRw502oOL62DwglVtfeTJALO1UTa/rCJ9GmhBjnZhHdB
WY0eD+Ok+MJ0kxrqfC5peN/dpYsOZF517qHHQAlD18RK4HFDvzpgUFAKIdKolzymVd3wprsyl0jU
tFseONgHNkkfAMJDmOBjpR6c/taRkIeAGpQvjfPvmI6hfXRhBzu8XSYQDP7ToLDsvXcqndPBk5mV
7vB5gK8EsSj9RijV3tnJ3XVvKXPQAF4AvoKy/fNs1rWmURZ1Q9RTi0NUc7BO6jhPnLnIGbdi9MkS
gcKgYSZY4R8ROa5kBLGYSQ/oFMq/+IkLz6lvMtwnr5dK3/ic5hvvXDISZ6xL/AVOugCdLU4vP9qs
K/eXxGQqhEocoCxdbKvLo/UufBByXuAGwNYcLIWPSgYba5XCPYaEFRZBrcSsvHhvIQY4pmgzevWo
5JgLvVJU21QzZMgqWt4EpWMImIt9pHGdLIBxa3/YVSQMPZV5Y+0THtle5fGlOhBmcuQUz3eJezlB
MI7uMG+cSTE/FAoWO9LeAfZdRdY276AJBn5FY44SILYGxdvsIb/AQkinJPkoQTFZCQVr666jaDOd
/Kl+3vEOFPmFMVDes/4GsEy+taw5Hey8zv7gUrNR3ZhSz88ZWblPiMePieMG6gusvRxLU0XTxl/D
i0Uos0w4mkNwo9Tj1BHAW+QE5PC4RapbvybHjT7X1wXTa+SzI3duWotbWcilIB7kWvssAWqv/xv6
aAFIJb5BSruSSep08aRtys6jlMMcWEX8iIKfIDZiK1owy0IVqoHqpe2E4oHN0SVVBImWjuU3ldVV
oWoY95GVtpnepyHPTdTzO7ExVs4IDmiHcBvaaVRu7tKOmyYtBr0R1NIkeBkCvCnLdq6VX+tSmezt
ijJDZRoXP3nZPuxt2sHW6lXXyZiBFj7vjxuiAoOYU/f4Rqj7ZvTxyeyQRHoRIWIaKEhOyBBIuCNS
HZN1v0r/jTmR+qVoheliA2Pu+kpeMw2q9W9ykriukdtwg2VYJtoNS46pd9KY101D7t6FAzEKYMKS
aAotQedM/Bharcf0o/zTR+OR5mGu4AA5VoTfbzqwrbgH9FhIJU3q6HsRacTkttEGf4DzXMee+/R2
mWHedajS6Z0mS9WNTfKNh0+cPTmKmpo8M8MCl0iAfiaK47GjAb1VPJTevkNOd2SxwF6WTiCUiQyo
HSHhB+jGm/QYm2qxGA54UfmpaN/kw4v43iqn0O+2hHSGMsb6o10RAiA/9D88m/EpXMarWGTRTDt2
pvZekNZbIiNwIGzNYuiGQpSFhmSgGG4Mk4oFnid0wcZImKcgXhUFVl1elCFB2lgOiyMQ4ic90uwj
UGh7kKzfsvgMabRj3IcxPmndfpHkIm+3ZOoPEh4qwqH/2z4qoxnIuI2pPjN0Am617NKxJcjgJ7dr
n0FB9TY6RIR08BZukRUV2WSVfbYTtlGdAYeQXCPMPJhiEkpLtirRSRezn1pq7d07xKS/QfDvDQaN
S0JaMTUsjyQOkLCC85BA1y7h39p97thCBe1uNc7gtXYITDEq4TynXn5HhxMhfZ4p2rnXGGNAeEMg
KyJ3LiFaB3QbHiH0EHKxOWi+TPEwtQpNYtSboqNsPYQiHxK2XExyyoKdTZAJhUTa9VHlAjaMIM4u
T5uvJxwuNdbdluMKh7QKmKylJLYtej9DRv5mQ8cfYpwcu9I4DdF9/RuufP4M8njuXiAhB2ftkuPO
5el0U0yQgxHhvYKf6zsUuUoTvGxWIHAWQO1GzyFgXKOFBLOj6HMIs1l80I8BobHpagQwFuAx9H4C
AQyMCWULKEkRMJdcjfg+tCmkCdEXUCialJOkrlfqVLiN0iuuiSXLElFqCBt2K7L1LOgjntT/5Ek9
BtwfabM6bmocbSYJ0R51x7ByE/1q50oSoE2/55r+ey0xM409Imr8Aj1T31m0CaWke06JgEGb+kSU
uY7F0HUffxMi2mrF/QS38HMT4+T3MV+yYSjBBDNvqc6mmr+eflNTu3uo6QnhK+m6j8o/z/erOtVH
l/y2ANMPWQOr3e4paN+ExZ4GNTHC0aAkZTvYRC8qir+zJ8jTnkN+rd3byDiYYKNlbuiEo/ywtB68
1oCEDP49E0XyewdmxAJIRol7HKHSmhkm1Umhfo6j3eEnECi0glgNNmSEmJCcLd9jNBopK7rN5L1i
nYr1+ZQVLv8RL0c5ZekyA/dP3RNtpluMid3PpaJcdNc/o1QYKUbBPzwVmVDph5tVG8iNljLnRM1f
r+Oay0+vugYwsSXhdf42mkbnxQXl61uolpOaPNGLZgJLygEEBG29jkENknGKNCUHq/5SDjkTXXT0
tOBaYhGeXP5a6QQX2T5fbGbMU72SEsdQcjbm4RjNvUXA5IJPUKJrIOJvpdMXJp6p5E1YXbRbbbsR
CAZNqQ3h2KAK1svpAO6d+jKNJR3W54OH9mzbdswW2xE8FCU29HfVcb/i+EjR2stBx/idmy3TwtvS
ufy0W8cpUwU6Jq0iOoBkLmNMOFTUSMUwOa8oENSwJ8JNhuhqRMl9M4JpNpArUVXUfIkn2QnhHnAP
PYAVOZJzzRnfFVR9u8WGVrToO6eC8VNcZR1p6PlJvALmhbWlH1D/hPw41hQs0oF6rqBsuUOWDHAw
wlHVmdCQknKJ0NpJp4LTCKxXRXjCRMs/MRdM3yU78QmgEJd80Zc1559rsY5YVINAERMGsYi5fT7g
vpC6uiKGNrH2xg+BfBYy+db0I8I6lslSxVB+FEQJ4Qhr10Qys2UA9Hym0EvNYpHkoiXA773amife
UrHGYIfZNgU1ywXmyaZ6y2kZwpIGnYq/a/ixGH/JOdExDyw7WgtUM+mCE6H8HQQ4XPnuCwc9mxyD
vZi4f8CAkmLcMjcpDdUTEIApqp70T7b3uUxruu4TrFVbpR7p/ISmlCai+FRZ8XH06ud60k40tEWh
LbLCPSBdBKVkSU6dFDUL6mBmaf8T2TREI/FGdy0d4asKi532/6FBN8DSSerIuMa6597lRVtZkjuH
whDEssnKvyaZQAIYgeQbe0yt0Ka9JrWhp2FIVyq7ac2O0HMa5YD+ike402iCUMRe1VLzUH3qlfWn
vIu5e4dgT9uvlnLu4yYFCB5xa6BRwGORiteyKPdbtSzFJvgB8UyNGUJk+p+2JPinRkx0REUkPB5d
D5p8SDsfq5woLI+LKeTZ+veoGrbzwSRf3ZxzyzFYVZWR5dZV09roNc7lkOJUgIHGXM3hZweoIO92
Dtb3OVwrIyeO40+ZrTKrKiJrCYv2Avmskuw6AIXXJKxCdavRlbJAijeHLfC0/4UgCjvOQwgxSQLV
+juBx6EBRbOjc7yN9ZMUo5/fNCfLhcuyxuxU+A30RngqcGVECVQ49Y4kCeXvaf42qR5i5NKIP9T0
NXNFLTJDuZr5QZRNfvvaSEige12MYEt0NPN5b8f6cClq5wswaD8LyIXHBv33A8uEooIF97h14TMm
SpU+aPENbdgdN4dvxw6QerYxJdhYEXPVCt0oEOuOB4qxpJ8OCoJHspwBjtJ6QG6H3bbZg+O6G4J6
MCbb1aQsE1cHEjslnEjfqE7WfGtIzqw/U8snEGIngn+6Clsp4DuoQiXcIup8CgKPg7d2VUcMDz43
HdC7/mAPuCClBnu8jdEs6s2VNKj4RKB7ZmacyKg8U9zS+T5++7maN+CFxNnjmz7ghhinypVB8+Ir
QsZuI3AjsG3ghTS09z39G6P5zmDCQx3snkA7Ra7R23iyVj9hFd8l66tRoxbBaDDItYOqxcVXeyXB
TIqAnehW7C5kybwF3XUESiTrbr2AMTdPdQov9YM1Xfxu32TjjkGzcVgH6MEqkfugSpRc7QBtBObH
MmZJ94hjwM+oDErfou0kMubhcOWE1MZdqG/LFC1FFHUL1QJRkq1KLykO+YYwiVgJxAyuZqHnSlC5
AoXPhRbIfkXpcX6bDn3SFpkJ/bFc1qAeXj/Xw55KftdO0QuDaVd0Cm4i8oxP7kxlNPsvqNBaRXJp
Thk6P9YlchrWPqpmesRtAlRV1UTKHa2KssakBneYWuB6YAR0UIHnNqEXyD8lERRyE+DfYjBrnDSl
/RJLlNG3lxSSL9T3bzSDQmnj071TV7bz6pC/NCTKxXEB9LynoABUoBVo8swawKBtC5y54OSQ+nxh
ntPe0xfwcVUvjKmeBne9U/YC/+KcZf+tqDOHsl7Zp0u2rMrjWmoOvj1UUer0OayTcgBCyUDxHiZp
wuUqg7C2zh238tn4wCBuuqBUuPlOjOVdba8txnA7exXcj/udMoYreAgiOKkHJ4sYw35+U7GWvryX
bhPEsvYzDN2uXWd6pHJKQFLbFQWxDNP8kLyRZk7SCbGD0d7zaSdgT1dVqlB02h5AlEJ3GrYJiylm
v/fuNstGihLEIwg0RqReJRkA+r5zi9CiJAhl0Ay137agwkpKPSFLd2OZZhR+HpKJsb+GgRhOle5S
SkU+aXPP9OTtX2/tY3lAgZW3blkHitBBLDWFVnVnAS+URUvv+4r6WsS8DYj5xrttEawF1iTA5ey/
pgrnv3qEXyxViW/yj7jVKguBh7QkT6trYDhh2qq2KVty3P9V/P5V97K/Y0+LdwbM+j/ysG2KtqPi
RbiKFB0rL+FuGOucDSbgCfLcNZqyUw790yTZzXyfWUzjxpzDynMEDDucOfZqsGl9BXBfN5xvFz3q
kMruvVQbljn61uLIYhpjAPdXigfSMV2hOJmi+6lGAczYGOQnodIvTrr38PLceWsgSfqPKCPi0ZwY
xdlGhcC9UJWH00zBHULNeqhuspm5uDAXP1k2iDolfMdqq8Nijrf+fiBfXfuQyfKrzHnnDdEOqfyS
ZSE/oCFSnyUl4IIUxSfK2rZc8VSXHAwL9G5BV1fUuDvgSKsKzvKOvMfPRwOmh3iMzN6fe4Xyb+S6
9db4HjZRuV6wF5ckswrMZZnySpdZ+nK/4Os/6h9LdymKoa+JmwXZx7XV61JQBFPzTP9ZcrCCY4Nl
pF50Ta9hcXGLf4Uy+POSZmzRsUINjUeVvb+CHT0/CK/iDTLFWpijaFb1BCz+z4inrYZnf5t7rgRU
9kuAO0YW3UanZ6bXOGN0q6wegk2JctD29P0TzHkVeJ1FREBaghB1PqDuuhemXnNS+HN9QQ2nMPdy
PdQ2wDFzamcScz6vQxvqlyGgsMuHy6O4lVCCLxVaWfOtWeVI6Kw6CNJg5bFRcepKCG2c8jKI28ZP
83SnhTOT0G3PBT+ZzMQFFF2xzfcflRy6OdzBq1E51RRt+9B3FygRYGOKeV/Y11k7YwSsyogZ/UPG
eG8Ysg9O99PpImnuEvmHdTqWBqh8cKLUceGw3ZYygo9FYruTlKV+L2tNcuRSnnvmmC4SSRmI4dp4
47T3Rp3OEcSxWY69U6citlzt//uqiaqKG0/Albkzb3/8l5Y1Y964NEzSIo2iNX+MVRl2rElX2Viw
sQO7ZP7qLVEVucm0mny3V3Pc4dvPxJsgcOu/yDsUoiOBCTrwFnrLA7lDmh4YkYDVXga57hQBg0F+
C/2BPcnhkJCRLClzhVaaBG09vtoTNxDqH3EfL9uST+RbrwEbdRNgJK7rwDZ4d6JAGirIx3/eq57C
qXZ2s6DUvSYd05hStppwXhV9rdTVyffGldH8XjglfBpD6DwohTLWzbGqEtIjeNkT1B44HLqhSyV+
L66BR5GjbrQi3i3n7IfFjcnGSx4Kj000owJyAlcXWcrp86hhhd7L8Mbad26MXWHCUXDqxd0rypS/
+QIPUxLqW1sICzxjLlhqQmEBoceg6MmiEAWpw7ZH50j+TMWPQeG6nD0ISYBnDgyHUMEje0HghD1P
1gm238Ni1UamkiNxZf0b8eO2hi/wGV5VXUlSuyOd9a001rc4350x5agfVM/iPxNlk7qXL5SzsnrF
vOjoavRHcad5atPH+s6+nqk+L5SQu1+WNXpzyQ6QKDlxPYTUUhlYiiSmofeqy6PO1ywlRilbbyS4
mzDY3h7IG7XOjMoAzZGGmsnJTWlPWOHNMIQE+ilFERwzVt/EovJgA9p1CWVXjSj+pSCIYI4PsR/v
qYmJU3wBX1+UgPhi9dzAWMrq5lB4MG3DaIn9Z7pLo102+LXIcHpHJNNVYUp0/rksgCekb0eQFkQ8
v9uuIRwLM62bemSA+e+EW35G+NC1BNqxKzLoJFbY/HIfqN9Dndj7bHGivECFXJH4UHVoxheXSVdJ
mnuV3S5z8UvMugRRZVVyPUAtm9tg0VPfnd9mm5ukST5alzSNo2Gn47gxbBp3b0EWTpB6IcQ2P9by
9ytdkElRxYt/PIYZD89uhwAc+AR6D8eKyqjTaOGcsIOTLiBf6zT75+5TyS0oN6T/KFTfjtoJeX6S
YHHTZ7rchzZ0o47NG7lat8EvAA/VUy+7lVE/ms6WRJZuiVAsOyw0zsdM+LdVO2YfGZEWqQ2JZaEZ
4/S3JNWm2V7gDRWiEArVeRqRxsEA5ylh2XUFoul5ThYdZaQj7MRFNPlpVaNQAmKU/hMDh74/AVHO
paZR4vE2wwDG5wVgHkEz7/YDYlVyDnE5FJLVWTuq08W03biMyU6L+gPqTIPvgKfCHHTxRyGYaDcB
kMNzAcFakRGK/SkeeJt4eXr+IBAslMtPPQO61FJdV3XVsFVyjBgLQq/fkHTM1VnSj6HwJrvpsLmx
jyqHSDZgKuq3v59ize7alpprCqVBMPnPjjUSh9EYa7jKOs2TmqonSt81WNX8ZHrxUsKr4NX79gHc
0QfCrRl1Y+gujRPLlPO+h8u/0U5cwLKXSu0oaw3T9U0L5VRZtX2N74XSuG8xdM2bCmTd1XfvorN+
qmJjsrE2VNMAzxJ7gs55XnPOx41Lzo04fxoNnaX9IGuDAqAi1gAddkJge18iTQFrqIuhnM8EmDRt
xl0bd8kxLNN4jZKIsdJTQqXRNbyFQMCdZsRaI4oAW5/NK65h4rLnS2ak8n0DqQlA2Dccjp+CzUF5
e4nwY+AjRSM29AppMFoU+EkyNGB0NFKpIBV6bDa95pz5WqScvQwaJ0p61NUszB236JlQHOjxXsSz
WICo5ZB2rtIDm0cmqb64X7D/mC0QQFqe894jP/J4KBJ9jAehQLnX5bNJQhxDZGn9tHngR3sVECBc
Ngf5b6ZQoQ/5NN81XeCeXJIlKvO+Rr8NNdQJREoz6307F7X1QrT3jtZGb3/jGPL04Q9nAtEwEJKW
G4s2jjuaIltSl2YtUdSLLCaw/qCWKVhlk01v0D7XDysuKdW+qD7nZqZRMW3jpzM39785CfjoVJut
cqPhLvgIXvr27SpDwa4K1qot4LrngzP0NgfJhuR1OZuKOGhsZ+dxxU+9Oj9hIuUZNeM5MT1ZkPbx
QKzd83Oc63IztIiTHVBUtZcweMNmZmcyIM7KZrcduFGRi6wCMZJhsC4fSmnZ0KXZzdt3R4wdDGdG
/nNxAhO2caxtVuUG/1eYruhqlz2k4QP2kvRTM/j52ulCHyM8j4naIGHQdWoOIt9sXKFmV/Xyc+24
traEhdnlUxYxZ3JKOSEBqSLxg7DYh7avybrnxwoedJ94NkoVmfOOfp7qYKKrlux62DVKQ1MdmL+/
Oc/ja3GMotRGgU+EYV8nC9feOuFSrgBp+IsQZ53KN59y7hLO4CExzoUNfiTY94e1gUNt+o+03kyV
DZapBJSbjdTTztyx3u7DkQAJ+VRGPbbnMLhLtDN4jDlPkf4zI2Gu394iz99fhNajfnU0Hd2leAyu
B9D2cD7cxXWev7SqX9nq7Z6V87li8qNRQwh1DJ3GJcg1RF32G4on8DB9DMaH1En3biAUSj3lFffS
aMHx731lTZ+UdvJI3nl0TGC59RMSdLZ0HWpWCLmdZ5huETRIYT0RTFo6+GRU2sb2yvNqlMiJR2/g
aXH/QHNXeq0TufYNWg/toEajX7N8CrfwPr5xD+SfG4L257UfTHbKuBbNdwczW3usz9B1T2+EZzeK
saLICMYtwFnIwWQ+rz4r1IRrotiJy4LaJ0XqRKvT+FJ+RlNk1t73VCWZH92IrxifRX9nlKZvZCz0
DGYAZbItnKRQQd1ZtNjJ2YL9Yb5ZtYrAy9aTP0+69GNE92252JBatCUEzCa6F4KPcgeaW2zMyR3b
Llsxgom24tUdYscKRwm4hC1qIZdLYa03HbZsfXYdZXQFuIMIiF0ZffvezxwNq6i8dYuFyDmCmONy
HdSZRIM+UEJ/mUPOA9qHw3KzA/9PrU9/JveRf90OHFUb0tlR2rRslClKw+GlcCoRRvcjLyeI0Rsu
X0qVNz1vP2UUYwCePCcZKzk+x8Ww903levEzhrRcEhmL0/9RIPk8BSTQprCxlIfdRQez931xAe1j
mLIkbFtWcxGS5Q5LNKcGr2Lk7X2k4pG0ZMeY849NCGcpSRdOQKuWsJdMpf/i/puUNc64bdd7i3rJ
wVFOIcglXujZhQ2xqeixXI5D9SRTz8JIyH7lFZX7edSPD/3x1LGd9L26SKQfIEi1R/gTm+5IdG5s
eNmPOnf/1XMlY6931iqwbY0J5lz4EdrASL0zpUbNs2OBUG0HvXjXmo4vAzjIcdRIN/mwKV1nq9R2
3TfVQ7HGWbVAFi5Q0JtyJGByz2GoWqvDvlVd2AUkcT9hUIS8XhSRg76BVmmva04x7sIznnPoOJMp
O3jzD3tPSdssEm2LEKyqDhNOXeqbUUFVnwIcTjYG3dk6ux/3oFD5UCs7vgqZ43LcffP8dBQph8tX
JbTrGXUj59l2hZZHogu/4YHLscNwAgJztMahco58v95awhWrT7ZZJXBjPlcIkzCBhDbaWsZCXhMs
N3MEzWJ8IFh99Pn3HKDZSXNTnbE66QhWHNaQGeDvwpbRjih41Ql9WcAsGqovrweDjr1qS+4XuS6b
CTfDWr6YrvQVKOfwdg1Q+u5sioi88ngqdYCvzbZMNaH5cIoMzHHU/8WNxPtlSQSiP8QTLK5Idkn/
ogq4t5tD/VrN5wpYU4mqFeeZpWsrDDsTobIoHDEpcZPdYo3yD96tNDIeSoJUpa9RkGH4cO2lPm2x
kFzz6ioecb1hrhy42EzdMaQt+qxQLWAk1tkPi0SmIHccwKJRd7evhRhqgKeiGXRpySpXLqVXxQuw
E2vY4qtXNUuvzQUYjwQX33hn4yNOcSc+BOh7w6Kr71Rz/3V4lZdXbHLfgrLF3i1F/uEEKvdJCGlt
aZxDTWKIwXTjU4VDsxHFvRNoYOrHFHwfuiFSl4pD1gzoijIDyCxbcXUw8lDdFhWwsGGOl+o9x1bJ
YJw6Hg3YkCud8OCdXLHvi8zly97oryVbwJAhrPm+2Wq5YHAH19e7unI/8oVSdnjooZU3uA5k9065
ffJm6Tr8qvwl5DKjqwH5MpoNmW1UCTMtYkKrRojK+0+L162QibS2eD+RDf0FXkRRmD+k8aN+VkKL
Tliy641lKYSRg+8uRHiNGjW2579+OplkXpZ4mfLDRwwfFzXT2Xq4WdjxrLgW4hDfOqWhhaFT2ZbN
L3V2wL5HFGU6H1LJn77HtceIBhR99p4mGKWOrWZM+cLVCTn9sjxa1etu3EzmW6lPnePc0ykEAkUX
7zB6uzEdFkDFpEwnyUlQcZsWNztLI0SwfW7uqiFGoTQqcxBbRpK8w+niHPBE83fOfWXpBxBisYHh
bCToYdfh1ZNsmfZntJ2Odq+OVMFH3VEk2v4Vd7MJZFd1/7WRkgh6Ne78zmGkZPQakvTkq2nhlIe5
np6IFeqMCWZJLnxwnk/ytVYdSDIcJNcRzDRMhHLerBdK9f4ETLjSLYWgqGPKdDaRm8E+7282oD4u
7pAK58vemmnUUZqTGNmnm5ZKNhE+Wn3yqD4NqilFRxV3p9kEjMReKTX3jZz6EMuZZaasba8e00s6
OZB8YVq8T3Gts6oQIty+Qh6NJneJGWoGVby0rY4/YmXvdKTM5veJN8YHjgi392BiTSl1cL0lvVHj
ElFVJ95J33hyoyuVCv5O3AlZIm6BsDMZ//wND6dgW283V8soZfZHN+w3kxWrmoXIW1AcMq5uv+iB
AVim0hcjNjntu1RijOc1Ku1I/jqw/1E997b+CqUUXdhoPuOSk5CbRqbzHCXxKQuG3oFlRWTEP/Vk
YFqTgiyabg29WIdaWxQLrDGw09mFLQDhns20FbJMysPc0zreYEA4U5jhtYBrS7QGEf01L9MRPeE0
coGDLn1wlbIdUFYI0AqyZ7n+TA+WMHyMWskc+PRRQlW+NWOCPibBqJLd6Mg7vE+xOjprCvpLNpCv
e7H4UBqtUi3BjYIf/VrRJ6sTNCju/G0/6anaxWUDj9SASAH2dYHdCW/SLqWIX/ANU+ABu5W6qV1L
8ztDWR6wrL8A2fliTuH3lfDAYY4ZAWk9NQ1iGSXECOqi5XhbEi875b3YaxdeJYoUmwRc6GEc6kJD
ffa32VJ409HO4V5c8fnm15Qj33slK6c5mKDxOVzmYOMnfff4CjS2N/4XZ4xW/HReVwAn0rNnfpkn
TsC3qbjJ5fk7gK9xpN/XJkDXA9mPo9xQCbfz4BwKkRSPLpGPQiELGyvAXhdlLFAcdCFQ8xjE6tZL
yqiY4okCnJMb0tk4Ons8Sh6Zebuah+x8jdOJ7xhRrKs+NMNdE/qgaDxahkon/dod5XoiGg0dk1d/
j5WXhI84PypW9Vi2z4DhEKALNf+nR/dX2eYFWMGyUrH7MkQelDxE+oElDkSE0SVW1ryg+alGqWK+
/lx9PhFyo1yL5/N5XLepq5qsbFXWOZ4jQ62I1G7LYN6DjeRwn7m2rP/bIac50kZf8a7U97M7I0Cd
TnKJEnjeue69kQima84thG6Ilzzxak+cxpHbRM7O8egyQuEi9Hg/APWwEj5Mohm0KDH8NDJ3YCFB
2Lauju7kVhF5dyWoGRR6DhyKpnETM7eKTPpzcROhgqw6O2oeqK2WFwkaNhRERu13cVuIQ9DrUs12
jaUAP3YszPs/8jHCHQJZCRnRyfAhuBbqbq0xEC3JLj3p1s5vh8EDaWKzhFZp09jc/UpbtSPMcuLV
i7wDly6nCy2kd7B2CRHyA9m9gd2mWgcVmzH02jGUJQFd+t1M5HDUiiel7uEactNI9iOGhaIAumwJ
nNpphk898B+HbhyjbeW1kNKtWMc/lvhan2Ksv+5GORqPXQG/mM+Pq5i6Hs0QQbYviwaOV2NicMOZ
c6AiuOOL9xcuu3GNxc5bgL1V6hGds2occjJNPGCB+Qzv6tjAfMn1YC1Wflj8XEP9yeMYXfmzzGQq
PNVFd6OUeamstAPbCsPLI9bb4tKyWjrDYOsVdR2s6sma1eyY+4hVJz/h1Ggj9D/8ET9tFsrjvfRo
/rN00VtPPp0rf/5PnJHCEZ1wI2o2GO0QLrgZIVjKe1HA+ohLjZ/Q3SA9bCdBzuEK+uI+b85IrnCm
wWRF6CQwQDyuSDxJCfAJldgCnhP5eV8ZGTRRbIVbye4RWjtjJGj1ziGZJx994w1YqIO7O4WxNabs
sxbI/GM5PDqOEK/L7NnUO937q0LaprppHAbB55BjfvyUA/nElrbpKKbdUsirg1n3ZtLle0Cmb3xx
cPADdzBtef0vKB+w8+lDWN06MRPlTEhr9OAqPav1iHxgANiMZRO/ayw42QStrzRTyMPkUheUdRVW
8M0Fee1dl9ZfyA1Q9X4RqdpKj082w8Zzld6QYSTZPCtTVsgceRTE/rIwvdzqcg4Mnbm4y2V4gkFx
Wb0iWi9R23TNKCDVl5GOHNP79hQEKjj0T95WtwDKbUuUNZ5QRhjhBwcj9p8Pmuum8sm4ctq5zpJU
Qfnu5IxOPZZ3BmufdXBmUFj0yIQ+7H2jSGpv+qqiR6TjuNK5gxf/BnOX/ARZGCBCr1rfpbhRkbME
mMOCreM/ELdyYC2aKLaY1UNHr0s3OyPsqfwGhR5z7ONsEb3K9Xiy7f72TP7Q+yClfqTu2DtFSdjO
Tki6b3x/852ZKgJI0ZI71ajx47JJD9tcMzPQAZ3JKvhZpyfWb2F7FZmwZSJIhDt281CKSjj/kqCK
h+1NQX3hw+pG2XnQGYgycCS/ClUXsDXNnz3TJSLSygjaeMiWubEk0cXA7EDEwLNfChqLcaFt75wu
MVBKkx1ULuxWQDWv8KgiDBW1+pykpkryY9jq0aLgmv/jHaMF2nUXA3YywBsTZRduEWqBehSHZgCE
/Sa9OZVPgpZ17lgSJmIcfPynBHxW8dyPDsalvld7zJgGU8f+zkNkVk+wCeYbChLJd7F2JW1Nnnng
mFnthyB4aw1vVMcZlXwY0WEzOGqFjqXHVLfkxjLwlZ2lAwTai89X8t7VCeUs+mOReOGlpgt/YXOm
lSYyvYG4OSQOfLusSvk9VIMz93toDwgduOEb2NNtj4tGdhkxwGf0N9+8mCXLiQgKCHxeqquNai5Y
TE+u+whvWhW4IKyJIatA0XFECFt6/EI5RWzleFMS18QbI/sK3pTCO10EWWiX0kIYO9xKnhCsFb5/
iFaa3fGKbKnBRSvZWzHhHT66EvPgtJWYE77SWkRq5JaNpqmoHepsr+xMyFW7pGxKY5OYpqM8xlwJ
oznkHAw+eV+IMBQeRaLRPxVbRHPWId+HALRFh0n5qVFLaoODtmiCSKVrTAj2UHRlJxBc5ofhOFlD
gtPKpEFyEcNv40cDlemFpkppoY4SGGbrELU6L9USZVaDYvoWGtBUiI9184QTx34mnT88XLOmWcSY
Cy1cYkgeA8VxVZ4xYMN4Ysq+Dcoz/sh1XSmGNJBhyeWy0MKn/AcxtCHT3yWrO2HFvjGEPSrUdT4y
42X3ZsPeVHr+85B5VYviWVV7UTOH5lGR2i29nvXj+SCuFf7jWw4XppGaPyjR2/8MXJ7m7BYIObyk
L9gcHN7cht4RaORzWZ2wlRNqpX4XTd4U+QjtQFW8iL/nMuO72Sb5dfCKrCCRGkJjttEC1bVdYyq/
2Elt1BsbbXh+drm910o0Gqi3uFmeivUDMOSc5mDMvXPuf1lfBPesQ4X7Pwma5aecp+8pyzWkfIwG
WrDsrvTDP9On3qGG27oM3jbwvrl57IR2+8/gnpWlGf/lD66NuKi48lcCG2jNgYSRgIa3gm123cHa
PCznLMxDwGWMKIZV3CcjI6NzFwdXyNa6nC9Tuh++960TtD7y8T3LRhylzQV8KQ7pTu2tQ9gXt/YB
zw8ifxyoxSJM8t6JvkxW9tjq6Su9gzGDZ0vMnBcamF+Ju1WonzRe+/0pZpGKBZWjA57pMRiCsSRD
NsttevrdtgAWvK5S0HCVQdYkTp7GA0Vo5GIR6MUsV3QgCpdjDLtFWhPLp5HwmK8WaVmtvqrIr0Fz
BPCeuKPU5ldTu1yyMQLZnzF72ZHZQduQPnxZNuHZkPoGmSh05RynW14+ZviaqP76G/q9dcGNYqyh
+XsuvXAzL0Rydh4XdcGYV61UlJEW8ZATrxsnqOnAEvx+bnSc5n2C9/lzTUA2tq9or2apoJUbcHdB
+ldyzt8dvzM4SW8Z1g91SfjugXzWQlIVB8/ewDyN1IebZZ4gkEO6F0ys6WsBaEJRLjpt5xf2w91N
nbDu+iKM6FLPmhsaWTGI2uzWt7VoBGOUSv52AOYXQS7OJlqUR8GJIsJF5VNhVRuV7G8UcXlaezyg
NFRQvkWrPFUwJEgsKjTqH2n/Q9KlEnsdTZjW/ik/4l+sYzduJb3FD+Pl+omasHWT5T0ainqoGzuw
iPWAWRTndNBJTwaRpL2E/J1CJvCLIZSR+oNIz+8p9Wpv1wvOPCutArfXaABummoHEfroqDf6Xjc2
rVgSjiJFnxtQxr9heooArJkAYodtAmhUy8d7uIWLml1HxoyxN8QqU613asR1+8rAunZkHPycwCnp
ZqnOMSh4h1AUdx+yz8lIP8VBWjgnRdopICu+fvIjATSYbS3xY6RRxiv0YiQvsdaQ2GuWTJIQjvjI
LfVhrx8Tc29nD7Prusq8AqYSLrYuadj4H7xWl3N5IyzRi6kxqgTDYroDFP7iaHHwOqBhxOATOODG
NLREtqV4ZJqqZOHvI2b6jEC5D5Y1UkqHju+Ja0sSRrbLZXOd1ZLp0tnlJyoM+FHl6T8yQT2zZBum
rJvBhbMpdZadDNnjN8xAg+hHgkwpIU2lXH24ipKp2L+kR6XRKml/TYmwIgLyQyvpAreFFkgOg3Xu
j3gxf9/lr+3e+zf+Cu6WeWAUcZ1iLubSBxJi3HPhG4lYWUDJOUfWHUAsDOTwvmpjoXwjBTa2s8bY
nqRJ7bZHMCtO2oZ32VzZYt/UyhQYtNLR97IfRYvEZ7QQkZMWov+1VymP9lUXx4Bo2bUMi8+uKDyb
2UgpxBC29OGFQ0ec4lbn6N6/rho1jkHbRMcWPGrcxIndumAPKwSfMHje9hv6/rsLuFi9bbU/O/6Y
PgvJakFV5NpbYS1ChJpigi6CTxCsJ8mJgLk/2uzJqhnzLJPnVXJoh+TwcTKEDBbBcQ3zcPI8FE1e
Q4VNj+G6Nm9Bw83idwLWKSqKP65e9QdutqakYx1fOsxPE9pqtfNC8/dkO2G/wMG1N4EwGknP8yKK
JbB3ZLPwaXp0TR9b/mnhGotyoFNFx9dZ4jNtWcJNnnnRVSK190zkV0qCXXmADFG6giUOL0uEAVI6
0o0R5xUbQDSUIsLqEqWdb3QOWx/XfwYqhzgfaOQe/q4HH2kYyo26D7MIAoYE8t7VEh7bEgZmiwpJ
GNXcxUTXp9ZSnXfEvKVAtQLc0V0R2p5ZhwRzN9O5MWtsD8OkaD4Mxr+d5e4fTL5LJO2jfIG9lXwk
+Ce95lfSSScxsQVXHiWtRbJfniNeAsLTv+Q1hGURQ+C6QS+elOLs73CNOoQ0+J7PyuedEO91oTvx
TQMBpPUgn9RcdT2vh2JmisfhBq6EFz4kqFewFFkAuPc2QpgRFprlsHRFrcRrseu3fASf9UeIfGEC
S5UcvFfk+vIhSEEvqAa9bUiFJFBlCWnU+ttzhxeevj871lPpBFWPJHt6D/HTtT53FHSMX5nwI/BZ
E3m/pXjhSfKfEX9faPg/5gGJIg7DVgkUpP6TB44RKHZvZ4N4Hr4q1Q9WEwmTV2or0QAC8eAWFHue
J7UStyCuQ/X2t4t6RNUBy/4sEfTaYBFMjLcsGEtJEKfhuVLgyIvvWZp4sVUYFRxT2Ty7fHT8IJQM
KuZ3Ghzv/so0VEEOlx4oiYy9UDdDTrUpDBLryiStHOGxeMh8zsRwDS4mScTtx2cfaL3BO48kTVWu
75QboPT2GjgVPLeYwkCLg3jW5jfT/v6asBbF6aTybbr/Mdh5S2eqkMgH4njIxEDdHBa4/vnJXT/F
LsEN7SZgEPDBq0LWHcqo9A/j7CN1UwL3r3iWDWgKCSzwxtj2HTVicS8HinGV8kasFB5GJm0rrw0D
AFrDkmeioqh7fkkJec9qyp2A+eqKb7Jr3Z9k75oLjHgd4PMOL1F4cf5+k3vAMdnaG1ExPuudP9Bd
oe3AH1ov+iFp/8gavkrz9/duU+n2LxAIpzGPv5AkjSB7HFGV7GV143GfJ2EKflLi5SjjqV+88R4q
g6z41qRoBqUAjGtgdVItL4n3TCDNZHCP/SU7+cMMY1X190XI6hYu+FHCne2Fe0QmWPdsl1qFucT/
V00GNBB9eK8Jbq3u2ALohXZyai2P2AA9xdA3ZHti4TjwNQanp+VpXNye4nzblu8yCRKLsw3RYTtQ
G0abWwem9A0dMKmDat9LxQSAP51TG6D06uY/UT31DKHGFEPdhYtF/gmXw2P/4VY8c5rqorzJDpq1
k7sEbJf96Ns1V3/J+RleGetY5xYGeA0V4d2WVsaru+tl2CRijT3xEcZsEZrpEfdfY+iTKi46lD9m
IkWIUkLE/KJUAVrOoeddSSMDm/0YSdRwC6xMjmiCqWo1aM+uxuAMzo42UHr2TrSD27R+1CCBFrNO
2g9XeAPpD0iQKzAb9sjOn36MnWT2VybY2BHUvl6+vSxelIikKsUeF7QYF+F1z/Se5GolhSB+e1Qw
qlcN0CampbNP8G4DRaBqMRognS3ZqqacXgvUDydJLJT2UNjwKdaHazp8iICIF9oAoXllNmNoNYp6
i5/SnCwylrwuYOnT76sH7IZynGMkkXnS0pdYxOPu2Ghef4jaGqlimMt7hkATjtyiC9yXTgv+AifU
Gkfu/4hrUVSTa0nsoJ/JTNmwWBxGoPm05XLvM+dXOH8Q8+i5bI2YsDz5/pyN7KFjScZpVCHCbeaF
CdYw28O6VUm9H18ekmWFAcIxnIinhf4mdDm7srFdFWxDLN8fXQrFcBHK+iRtmP9bMCzbMtaoNzox
oYd5W7JIH/wgDWc1EaeM8hpHYHV907dfPetDcaTd/PIID26ZxYWgkiYVwzZcwcRyL90N9c+I577B
hJ4aKcyEj2P5nI4iGFCXRZ3ckyTQjQHrwKog+dEBh4UzsBGzeA+jd6kn8GzvONciiGTQODIpwM38
q3W8CGmiztPGLfHzQHSfG8yRCkxAm4qDXZeGpNdk79uQqNzX4ye178PBlu1mo0KXGzxqAVqAudMB
1/2/wTDuUeEUMOliNqR3HNIruTV5Ubd0WRRZETj1Vu6i2jVCAjw16IBgWd/GYYmzz2vkaD0M4j+3
sOg+lVl3v8IHZ660upfhRzPGecglWeAlpCZE+NYAMBMp8w7u8riWZ9HmAdTCd44OhLzasprw0w/K
Im7ctEYZ/kwSeyej9IfgfSXDhADN6SAkL8XNwJ9jh5Dw9PKdpfIsW0/sAYxekHbm+k0YDBtEbZQM
Z2YSJIzFrRNt9puNkV4sAheZyHOuNmAwqYlMasUX1yxu63eX10tWNQfJ5/+0G5b2t1A8L/D/r/t6
CRqrB4zgTPMXvidZFDVcJff9hkUbV4W5JAriEs/m16yoxdd434hKYPK4RK16bHEyKHt82cR8votD
sl7gRwIqH3RoXBHXcIzcNijmUtwhgZS43oRwG+A0OWPjQURFQkOF6soGS7ywKrsBnDDi8rYyVvOh
QaXTFvyC30/19Qh+XKQz2WPQJjSKbb0AvLtfAC9VWuZv4hVSZ+XBHfHvTYXs8hf70ie+VYhf6eqO
Lo/7st257vVNAe1Y2mW2EXLJQC0OnKQcZJoRhXNOjKCI3G2tRfsB7cY5N7HW5Hgbycg3ZSlzkaPX
FVY1rFKtGynYGnTkmmj/2KjiNOS7pMmY4Tr3QcqWPz6f/0eBs8X+hB+FaM1dl8Y8ET7NMy1eht90
TSnOm4dm4dU8UTedWsIoApUDGgUpqydnUt+VmtoVk3ME2XOPUz7jYVvz1v4+IIJJ4+Gb9GnV0eO4
hVnv/pUswJWqdOMgTd3VIdnIYmKsARB/Q3fXE1GQ6NhLAWqjdGGb9Mh7p5pP2pszeWsmCWEtJw0Z
ym3FI/O3UBHGnAFwxNC/dyhYAggp1VxElheY8b8kWfg1R5aWS8RJj8JWHHD0A7QfGTHMLXYUNhZz
CcxY3S/D2B9nVjhFrl3ee+wEL/3ATMVW416+zTK+0G7lsdMMA9ZOM3PrIXJr2hdSjaJYvW1nRiqg
BX5lXdeE010hfAUVg+ISZNDMjPGBlj2Kc5EdXyyUnab+/GM8kimgGpZ7vH70+ksgUxEnPeg2Sj7l
pPkZGBfRLlUtaryOcbXU38WdmgAdY8QuvJKQUoSDUm4wTzoNPobjAdQkfNIhIUsNQGY94mLGJqef
1T2dOdMQODX/VnW6gBadaNbJ3QVeF9gDfqcPPLNO69b/gSBmOrnmTi/6KTOmtBIKe9hQO5JbbW8m
XnKFWtd65j+qcfLxylNR3MI8gV8kai4eTOJoNQ1LaAXnoCTjhcy3hGwJjLNOyZJ0xhDdwMuqky0Y
xDpISYylRTGPLV3OatP3z55YH3gR8MC9abWcgpFkSuqtaesxBJuhjI704PcejoQIN/BTTAd2dm7/
bVYRJ6qsg9aQX7JnALumJym0OrapMAmvHWHHvCp9t0kD8kya5nV1kmuRsO1ur5MQgCVxQ7rj8iQg
VWJTqDubm39xq9Nyp9H6lIxjaaNxXFU7POLxL8MnBT61ZWl+3n1PuXYgaNW/fqjyd6dDVMGKrDK9
oFCkqFOj6MSP9axV55Z6+1Mt6R3cDs9Rw/R4enKc1uHT4+dhkNyuiiYcRszDLUMBLV6XIoCFZA0j
1ZWuCHj9SXj8cyBUE17pwy1GLT5+uiYpmNjvvawtN8ama2sEnDzV9bFj+jxPglI4X4cHyw1PMhSD
BW458CmDL387/RJx3tx8Tchwbwn3m1uuewoSr/0ctAxZ9+XMHst8J8XwVnRp4KU6I7jLucJRqR4S
iQYdJgdbTG23Xep1ou53kA7UWLqsXV/GU4OQhbQZNEowJj9rFCjxYee6BCTABAdF1i8sF2hgWf8m
x9nDSyAgW4ilEvKcQKXmi+LVgP/iIK3AW2OE4WEgvLlTdp6nRdYof5sdgjSAFS31kfX8R1mc8Q9r
fyjfrLcSbZITxsjJqZAceYcBjrX+yRmQu8fDg8h23d/5YsKathDG+/PlMxqPS6aKx4MXxeFMf772
ITWVhPcJprHSgfmcQNlmZJUvQw+UubloQgJCC8+TCdpTv8D7ddaX4ZXqOTkZyXCoYhL5b2gmNBG2
N3Lt7mxv+FffvOH5Nrz1anSP5lqFw0NjsLSss8sXut6rdQsu8TSoKho5XJ8fS8XeQqFq2iNhrYBS
M+3Tgb8HIM3kvFd1hql+/+d3VpTj2zBP+fuhaeAAZyYyuMeXrSjsguo3tGg3/z2iRL8eIwWIOFNN
pJhEfx1dry9dio+5i2FZEY7ZOABd1LHbgwRpVkDBn7nIhT95A2zjnjIgjJCDAMHf9C5+DW23Zy7n
VkXh7Q8AL+ACJmtGkDYDJrXesXqGAaFNcfmgSr6T+qjoSIv3Q2P75toCHFQAcyI2vFj+P7pkM3ah
kNeOTB0mMP/19ArTEKuzRVGcJ0cmlCvJ/YNSncMMguSKd4j/84u4oPxmbC4C6aNbAkr8aasL+b0m
IxEhYFqzQPo4JG+O7uxNzFPBVHqwApAtsh8ywkgmNeQ92CkwQhwdjOj4eq8xmo5X1j8cUeLsWyx4
JbkwsYkJgRt6/WXM9dxJ/Yp/i0Mj9NKpiO1I4CQ3PlBqLGTQzTnUyNjLZlJnILovqSGDDUgjD65e
ye+kCzRFwkkXPN94rUM0IjOkhQJq0PzVn2+/W+tExMCa+P7TAUjOyRjpH9AxZqCXJnRGz8bEMDMa
PDlLrv+Gd31VwJrvBKJVs+xo12bY5PiIkeS26LcWIxp56w+eKHyKu7IWfuAeCOAmnCbVfs9+3a5m
OmC4/2qDpjy5+igLpfLl0f0J7wIVjKGheVXXRYv8OVZJdF3Hbl/+qIqwMa0NQuSf4LJBP5DUoiB5
O7QNhabRFZM8qhCuTLRghxk/juKrAxrWsJvRHjjFNpBMFw7RL/79GH5bxbpjMVdySPg5oIbz5c1O
BBDK9qZ2/4iJ/unwqM4x4mEM8Vee06smOQCZfky3RbMAKAAe7r6/8LN5HOVuXjdQzb8MgQ+5jLO2
+RvaXqtTPyY1glwpfzopTS9GANR85W6MCC7huBsfKUR4CTtPajgo9dxfiDZ04fCjthw182GGQfJx
wl68rJtss4BUF6KaOPVqfzAPDJudPAma2y7FQJA600jFxcjwFA3CVwkWsWKn+wN345kAxUFPIi1F
SqXTOsJP7wSALnTVcvDTsAlgnNYCeGM0Kvv/nMywGQt0dX59/cZS+q2slsBYxwndF4+XB7mypH85
0GLjaca6zuv0MrcTayScvxFfT2+mOUqBhWzVcPfOLQ+RywSJF1Q0zdPecQGgXwFMV+cZJ3OAXv/P
nHoThyLdRRuc5U+BMnDNQDwnn8J87YDHF+eisqi2mdlYaWgVOjwCfyYqY9tYP3jDxa7UL1HDD4Zg
HrwakX4Hozb5rmsQhW9PXP5yLIeMTzLQo19jNv61BSwF8ZGcVfg7DtY3Pi+fBvIxFBOj4QGo9ovv
Wr7oKhox+q/SWZkv+XU1AXhgamvJbbRwIvyMfb3wd9rlwoq0NMaTewOAzR/hmAYLqb23CNXB6q3E
U+r96MyJcSwPqQxFaw+47qTP8xWF/8lLh3mmPBnM8uGneX5zlMwn3dAJnt4+dmQjNdzf9xcuAgkY
8MHs5VDmO0oJDXg/ZI2Y1BmA+Xk1PbpKRbiuddTLtCz+oWv9idWFTaFnDNWUKet5kveoZP9c99il
nt6Qgcq737/GsAjVg+9ocQnc4lzxR1+QNiqBuNbRtmavgfPe4HGX9crGpjBYaJ4ziGN8GZEaPAVa
y0XVNZ6OXq8hBHCOwRTErX4d/thqpc1FjLJCmq2RFjvz/Sovpxk//6iFZwOrg6h6gOnaULggKwCY
ewrmqBHlciI3v69crMjqIenRCi/BccY/a6U/mLzG8CsOLsKXyfCLXqiXFVQbS+vgrcvVvijBLa61
vGB5aGtINx38aVDRMn2bcNzb2yopo8xTPizSMCWPAa7ESUI8ZOH+DcEiQwMTrPhTGxctIRTTeiBN
sqvB2zcK+XYrvUbCb8aAhCgHKB122ANL00J0N4KhzFk0n/yEq3ftAsUMfIYqlRcfZ09zwrV48WRx
2xPVaJx/iauQ3J/nhPF8tN9O7EfOSwfTbjWC8rQZ25KjAKVS7nPYzXI+br0aIhxA3Xt3R29rVp9b
2YSuIyI6+74RCYdyseGP75Hc3MUb7MecL6MIou0YUmbfRxKn1T6Nq+M8ywG++gq7scZL0QbsZa0q
PbPr3y59Gb5RlDkw2kYD+AeeGUxcWrpcBYMvaFZV8XtVmrYhGwGGYaRGTbgZNY7J4qXD2eyxhUMN
BBzo4NLLuPtpFh44fYlo+C1uOJc5Vwg8ykZ0qgskIL4hbkD0vX8AKdjCfRH6o3aO9qesN93mjGpm
QIPq7VYjct9Wun51hmOLl9HWsoRmcEY1yJh5tW1KniP5EUrf5DuoJ2T8H6t8ntaz7WjLhxSxWZpo
0TCCsA0+18SNxhQ8GBFBbnTVoLESnBKaE0vw2m/bOGSsTlNQilGq5CMFhB3LhrFRxmHd2ZpKIqh4
aa+nPMFgEjuf/lZaH9AeRbry6nEIdk5/uMPYAZvnZt5hFLsfckQ1aHhbdNqTs86IX90b9TNvE10Q
u89QQYSuHTcght9ePM9+lIv6KqP7w7gBIfyByV1+R3z0BjtrbR3eL0wIc3bUe154v7GFse5BQGIQ
Z0RtniT9nBZP1EMGIFhneN4pFPMiyQewbGV4t+of3hfuFdO7nwSLQw47OpXLWr9Sb+6hjyWqzSgS
oYQ1PMpCikjw91s8KAx47m3viaQhfo+b47TLwuDwbukmrOLHMxv+w79jhva9FhWO91kerYU9IYG+
37EExv0gY9Laeb/35dDqbP64VwkpsowsVNVPzP6v0IXjjBNbeg1J8wudx0f2q/JoyJ8SwlHqd3PV
4nSGJmU6lMagXulIc2olWN6abOIBDSonnn5ZFgpyVIaRIwQVdE9Sfc4ydzfwrv5W8kCDY21IAcrr
cN5TvisQiEXteSD8RHusDJ3R5ML9GuibHNkptxUAh1MUFzEWEEW8JH3qaG2x1Qg6w4rzYcGyPUH9
XimYm6SKwXec50DCF6oPYa0Wv5IvNfXp51af4XmOKg0YKuOKI7O/QB98Q3ZAQW2n5+R3TWF02FXG
JVEjJCuWQ2FucAbgIRc3LMwPGs6B35SrZPcY8+g4Gd9Egu7m+2HVf0iv7YYz63iY7CkIPE6ev71h
MsG2HAr5KpNfrE/buI+E67fORKfnDOxOrX+U9F5L2jhQ7M42pAcPjKIeVpmHaDDIrY6JiKqrUyeW
7H2sH7HPg/CK1NoGulgqqRtoXX27bhbGYHS8R8Ji/nf3K2yyo6hXYY0Le21PlJU5+1Miu+IqJ76s
6WWUw/R9PUEcpPyfeWOIRahkEmk2eySf/bgEUCPudewBClOD/zDBRvn7vlY8Ei3eD1UN0DnhA5me
3uNUhyhFSp3iDGHmWBfC5h0UyRO3mqeccrbvdc8CnYSwYwMrg88Ht1+ZHv16SDX/2vH1jEU0Tq6V
6FxU4C6XTyv3bLRad0ZveAepwNsymP1qZZDSoq845QENTsOoL1NQLX4B0aKx7DM4m74HH3o9Xe85
4u11p+thuzkGAR6HzEAczibToNsbiw9cvfik9P96pnPbO+xmxZ7qYsChNESt+VJxg3D0v8xDsDkd
Y4hOyw249K+ObIBWxBo2WVw76ASdj+q355/FxNABu4zBaaA/fjccGa59vE9bU0xyy4JL6nkN3y4d
PaNmvlVUrpIilrvpaH2M7cqA43zWYCIX3U8L466p4kKGVaHfEPm+4XPNA28T2+Y0kQ8lCsfdQ5eR
Z3ZaqEPWTHoTHeQ8aur65p/JGXQEjYABXqTy4WBnibnfpkNk5rZRI1Sczjv9Sy8vzri6QVDCFO11
BJx7u4EbCXGH2txaigDAn0iqLqrkGtTiINQHDQMpIc5KMJtiJQSi6y2m/KY6cIdG+SQ7ocgCufr+
kYcDNniTBuYr1LQoLY1cACpFAk8J/0Yp+3mvQUsjk5alrIen7C7CyWGSNbzVANFvZb1MvwNE5YpC
ukQqo+g6yKmEdkFk0QQOObbtLVg4yKPGkYx1jTlPsvW3QKD366ovQZX2ibuysapv0kRKawo6CPF/
uwTvYgmfxOYl5n2GurhDY9lp7J9krz66LUj3ZKnZvzI7NeWxPX681DPLGX+PsKDE3LQpdQRTvYQI
oQ6f7kpElvB2wqbBHbNMZZUBYt78QKOAg3MZdshSg+bwwAl4bC5VV+bEJTaqo5Vig6MnLVPvVpAr
UMcmzyGnTjF+uOf+vzTuHqJsIzNcHWcPAfLZZNFtDorHWXVWlbGwEbooZWkAUgMtcXjuXN6tyES7
sN8CA68a83lqGZgocAluvS33e1UprVkrjfXXaIdkapzUlikJiN+nwIpAXJBD9l0qU/DcHSuKrzha
vD0UPbfN+ng0SBpZQQXsS+MVTVZpGEhAlqfbTFml0/h8OiB+bNfMvX0kjTgTvEp50HcS1ETzWaGV
YKFZjAfpz4BvOJnkYgvr6Kpav6QqPnoHrKJLNLYt5AaDXxN1jvz8eFVuQPKZAEBBCYKdFVt2pYGI
6/diCCWNfUy9Dth4sRJJLccLlKAwouM69Jux7jN2aKalK7RS95ibRxy3cUdekiMinNIzhM4CZyrc
O2i8jMg+tVCUo1pPLAqdzqlzFtcJ2m9YPZXYEI1MExEvtl0QzupV/YyvW6S0F+PmNEozVPbJyqny
7MS0N1+6BfO5GMo8bD9/E0bvTLVWTMhjkuVpQ5pyWBrkOOCZKO4bBCGyy6hLkde2lKGMf2UHjxP2
nWV/QNNfalvzZRjSRT8ff/yuZcyGNvZymGjkjLV95Y/K/oMkb3Ek+tM84Vm2STC6BdfYgnn5Rhw4
EN7VC0XbNOAfCU4/Zm4ZF7bTkzmmULZNWCaYBnRu9oOjwyCMDbJ97CYnEivACvhkmcNdflskIQP4
OdLP3Jzkihp6sOsd439ZRpASX56A3BkpwzlJccQWQ7pPr7HUY1IWRq1fSliE7/TKyYQ+51diLm75
TO2TjPXYfKlesATlluBfaAqtGM6rZwTWVKbLzom7sreFMmwhwYhb8Ji5yo1/ahhhoxV/f7japt4v
lc7QgbX4FtRLj5lkYebBF83ATC3jOSKoheA7Le5o1Q3syVn5IJE+USPrMPu5T42SMsAd7RFDTmjb
gAiGlQGYG5Q4b9axLX6CGfe1at9N2DKjvihHoTWPawtvK94MWnEE07F+f95xoiOZlwoQPIHgoXQo
SqrR5pB8q4NDCmOvPmXUnq3x8AZskahJPTPMn4fovHtgc2bVfxOJogjAOCVnhn3fl5XCNp4SpRd8
D4Pcpz/pXYcqdnFKSzvwm92mblehEmKLqPjLHkTqFeJ05sKhrWFzafswnQY/pyU7ZZ618QyeCzUU
LGZgZ3vXy0tHRRIN+g38IIfNF+fGVUZhEvU6ViqGzUGwgVbXuLJdF8+DMMSMlbhUjYRnOzsygdOs
XN2jseAu5CMDBbqlQ95TCRz9ZWQAYw5en0VVdVN/CgJfaBxpJVnn52MjE0qBkQOQD1iLR/pnpSVH
vRmugweKu7c2GSK5IIHjkSfio6e9owrQKbrs5ZiIxbAVfInHZz0l6poHqa5rC+xvBu/xoHkjJCNy
WfO1SD+gw3KWH71kLwNRXi0KUrnnZhwdEJ3y+ggrAtHYYUb1zlwvrx7SqlAOEhgvE+KuuqDJwj59
/vv/lboQm79E2SR4iuJgawWNTqDqQg299F2XHBhxBeYhghbF4OThuD7vy55KCAnTo89kR0zWAF95
j5w1YxkbhU2196LEM/0/lHl5ckiaNrSDftA5nl+UyExKJIK/F5ODx+xUIBVEq3OsfkkE6ww9bmnE
yrrGDO7pgbh9i/H3Q6XtigvnYO4uZ1ttX3TMzh/A/0e9cW0VTNFEo4NwSo+afQRp6QypEs4NR3zo
YmTJfsbhE8JR3KGUSi7bKmvRsJdDOA2IU6Nb1ydm7KTzyteYpktvHluHpyg8JNPAOxPzWFQVuTlO
eexyWKZoTUISFDhjs61FOJsot4IjfZCPjWfO5LpGvPh/JnPcvuyBZ52IRY8s2EhQk0TT61Wposbp
T8OuqZEdqmsuWlWxJ+5RxONBWGMczig6zAAHTtsDbbh8+BF2O/UHin2EgdVj/QPw5eOpqJH0Ec9e
blV4jeWKLDKPvcsG4zxDqYQTzXvwuGJva6nV8RWtkWCIIkv0mpT//58wgI72QkrgiSW++0aVbuCN
kdGayBKxkNAcUqyc7JEzm09qL/jF3BisRojxTpB7Z8zPbSSDpIMyIzwtTl03SxdCkfJwfUDQXBqg
nk7N02sbGd26My5OUURRyr5XNpehnDcQ+WFJLZwapJyMTv/N4ht4l+5K18cNK+ygKUBPmTFW96D8
uAJ36NQkOKEHHUR3ljmjIjSktYocDjJYULvPs4gTtES8+PxzG2hYXmakJPwr+v/yxNMglJlIXds3
Nsw9pwXzHCGwVbSQ4TOnVvPdosNfGphWnq2xuhSXiZY3VY4yPprD+mM8QIzb8UdZOtvR6FWHKZ6/
3sFRCyDGDirVHCUUXoytyzZnuYP+mckQLfrVeC8VVyejCmYnBuX7sSsu0YQMl88ENanozywuc8Y6
bdr9e1kybT3udL1FlIYR/v+vmW4zER1VYXDZ1jBOjwOKpSxiEeyWsRdPd5XOLhf5wQHozK9N8Fte
Vwb1XDBENKj+QgILC1r3XXEXA5FH4bTg7DGXtsnASG0sP3ScQLCnBkmQte91vfwKTX/yrqsW2r7i
s5cmUDjVk75uKKLTxhuJhHvzKPLY+E0E3Bf6uWK6TjrcY4qGDOIaFT5wqXP7+S6bPlqAuPQtECNr
3sTQ0nmnHvFjn1pJHRwyszlrdMTd86p59D2Wek9EcYipSZAwp9mNPnpjilcEneafVtvS3P5DIdWg
xDCxN5RwMD3hN3HoVNt3fGHo+NZIslQc+XZFh7V4Z2XK5jnO6pG8ohHXApwB/ntXEIFiMq6cXKYB
SoyjidENLA4RSBTTUnJS/pZinVDX997XP1Rw6oxN+3HpSiGTRX7Ibbj6rBdEcSqWzIskts/+P8ZY
RUYZY6Boj+DErR7iYw4XxQelnGFJAnFZi+hIEcX0wTjxu6Gfyp5hvXdmJTnObnW5P/ostNwY1i++
gVvCuAgN92gOuAP44Dy6L3ttoqdqgkjZ2GdUUc6p2qBkUzXz1z5ZTiEhbyj+URfCpZqI+40H7n1C
MFTnjHmV1PeW8/tDy56PHlkx2Uop8lAMf4+2t++MRqj+dKweSKB8yfF5FF8o6zaR8S+XAqBGjFbI
7UeO2C/thr7R+nidJ8Hj5IiZv0vgNCJu8jXUDZ0GutcE/sHOB+mW/RftRb9Hgy8hS0WLYGjzLdTi
/rFLad1Ef6u0eClabfFVjvEFDBYhcvdvXEsT5anmnC3CbJR3mkrMLs8/w5Ei5bIrTOzIYi+k8SHu
fDR0OCQlESN7a7NQT1n4CVIfjZ08XYWOeL+2ifvIKUMSJ8HHmNXt+aH3FL+25BYgyQSq+ArZg9RB
Ku8VWWyeyeriMGpQkx5L3+QsF2WnhzwhwfS2s41HH/AgCOvoJW+KTPBV1aMycfIdR4Mg9vw/MMoY
1d4LxB+0OTX4aL58oLgP52szF1NU10W0lT4bC2S1M5fGiuh9BklEtMq+8kyZXwrWSUHu39BpYnAs
mOSShz/tYGomD8Tf2t1fkw4T3gKZtBJw8bme2fu6ywA+0TqR4shD/fjUE2pyDZQZ4GMw9dbvf/n3
0BVzy3Timt20GEZwshe7bDPvyCOL2oYVvcTIXtXlRclA8QVKlL8fSLfJ6fmXMb/xWqJhTSWNvGub
QKxxG7fS9QYRHQwgcWLSyc1Y+RCPsYKGdQ9lJARo8vs7HHcO88ps59VFBz8de7o6LtObtlDu9tAT
KlTDZ/52vbJNw+9bgTroLk1yr2G7vcuSlbhGaoIfHIFApNJVopIXPCOvuIH8K1xl+HaYlLuWmA/V
GaVJ3ZbhLBRVfS9PFEyvFOW71XzauAOXwk/dThyuT7WHO8wFOhld8mc9zYNFHg7QrgSO8Arx7Rve
JAEFXRKieXatcIp9KFyD1RXTu6+cg+J64b41hSBJRH6gYAWM66Wl10Mu5yJ3Jy/I1ShP78DofNDt
x3VZqckIXY1/sXUQXvTR6otp0eU7BDaPuF+QraEdyjBBIdQwA1bWFcStOwM/dXmRkI2eaKa4PLai
vyD3uSPr8x4F73Qw7QwbckNoE9jcfdMwlpKfmmD0ZzFrg6zQULvKNNn7NgrmsmjNj7bDLf5QdkUc
9mZN7tPu0Mq41JcP/82buN2Atz92+XmYWDCrxidQXbg3OM/3xg/W12z/FLFg8OYBfNcbfR0E3oPw
2RsAOR3uHCP3W7pYZS4dX3LN3SU1V7JC2/zY2X7n/DkqrhmiFvo+yAmOfKiEdzAIp5f3zKo6uYcJ
/KZ+GxzOOw1BBzXRdYpbdoMmAT79ND9Uthu6g04H1XDsXmSezMcOPgh1atk0p31UkLxZTziWrk2B
v6xrO/BT/yS2TnXESDXTuTaR4PNy0vW72m+irRSVWhnClNm7W+m80fhmK72V1lj21imr+35Czq4g
0/DfVIa9PkDqrCq44eYC67Bmo+K33lk9EWDjuFnBirtmgLUAgPV93zYEMkT+6c6zt++1Ehzh4WFy
lkAAiBVd11RZDHHzOUx5iXzORUDeqDIfaTITb290rGfH6EnBJTiQG9h+t2vJX5JvAT9OA9eMqKpH
vEgFoDSWlEKQNdopmjFkSf5AN6x5qXLbRKiVRcgpGSd/8NqAwB6EvfKZgDOt+JnJv/E0o4tRMJTc
oIej5mP/XDZrjk3wo6iVAyfT/2QbYW/Yu7Fbz3A5KBsm1a2nHh3sveeTnKy928rWw3nW0tVQbsH1
hSK67zPnLSMVdti0zJGO+sHv/u6onNezmW/Of0bQ1jx3j4rfOPEoAROkAaBJxGAfcG3kw6yMJNqV
ce3G1XECaiACTrqRd6srYuZMu32qsRsoDkNJTM8wri5PhS9LNcpsVkCjIjgoALi9FL7Q5FzDIiHN
b3KL95/3XbQ0aUGyxdk/dECXQ5Z2FYlRIRYUukKHtyDgTToL3mXexaTRgL3AvUSE8SJ2FpEr6imm
abgvChCirz5Eboa0uTfvifzLsrq5b0Csxvf1Ojo5B8pE9x25DvOQNPKmL9P9rPJD7asXkZ8hBFmz
xqo+TIjTf/B+iD/L7JcTrg07nOMXb0hFUAwd9+iGZYG+ic4bmOSKC9oJl1GGl6qfcmPNNGIzlRfZ
eKGL0q7R3Eu/gg/tFUFC4eVKYvTEIWnPpci/3sD19WRF0qFHr5iVuteS4KEUsJiBddIcsnBarMXc
Hk27t3UuHT9aDZtrg15BgSxsBVY9JxVTR5Hxm/fyoyO1m6+3+mhAFIwTjeBaB7m90wnjmcryVE8q
sr0VoZeqkbi2UdarG6V92sAa5G7dFPxnSJIYhAGn4Pp9w5AcAHbE6RuNMBhonVrV0PMQOg8RdXqc
IDdeqLXoTIEtFe7oiQT5Gyck4t3ns+FUu2p/X+XDvZAMCrYGpnmo3bi1w8zV6lOZou097V5cwlMw
o9v7v1r6duDqW7eVAzKUHJWu0ba2JbUOBtUvp0aU2sNRpKrtl/kcLX/B+iWvIbbcIKmVBsCz97jD
8ZGx7zce7/kjoxfrAQQ4qYQXh+UwnIp3bqj8s34GSdjqlXJW1syKmb8+1JVeImtJqsY1o29VqGz4
qdn714RFmpZZXHSMi3iBd8Qb0pV20wK6ifCZjliNEREqblYjG1LFgepKXMIK7kN/lNbcGsmkSE0K
GUWX4CbEpxJdZqy7dErq24PRuSCU2V5SNDeUBh0cuSBqXtbx2fqV2JKT9YXncBZuNmL8cma4X09S
HNi/RYuaUpk/cMuj2QIC4BnSxT3OqCqLzawadm0tuV6coZ0GhbdqkMsQUsAxzgrTD4EmmxDm6TWm
iLuTTIkiowHeCvDQGG4oJuyBR9J3+/IAO/1F9kcc5+SlAoHkXtqEyyIkMBpA+Y8yUl7LY0rCUJQC
gGLcgU+G4y2EjcdutouP4tQGUtaORcYrKVu5q+RxiXrCkpNxmKWap9eEh+IOXJIGwCBqc7OLgwpz
DMYjeasCd1gxJjraiL0/Rvl0r4K69CqIriS316/pYJVWXZdYH3DkN9+IksoMlDMmy/zXe1kZ8QwQ
HssEIsXwHu9nr4vLXn04h6ru3Ns42eMKvLUFSbZ0mrSwR6Ly94eMcMjQfOMyLPr/wiA+/q9h6Hj+
NxJrrXJSJ7ipD4GsTrWB1sZkKd02QDVVgzgcyD9jXUWUWpQgnI9tRoqTLMJhIZ5DIFG+XKRztSpB
prN2JFM8QjTuWjuRyDFKTtAwgrY51RXr05HwGzHLnCe6tG0YyT6X9oIC3dynluMPJik57gWqpbIR
eQni9q99O3WvT+w8fxIr8Bv5TWyV/2+oLDtXS3SkBYOEeecv4k342fXwVyOskVc+ckDv0qR41ptw
F5gepPbjSD0JZAnzXDWXw5vRBCscA2+uFAo1eIYtkaXzbCQMQyMwN+6W1YDs+CAJ5N5OiaRroAqH
vxPqWQncBLkxOlGcQ7YfIhnL9GXWgLzUIm7HZjWMmvlZ8uoBp8tmPrI3nm3o4/ZqWXrodMDepUdw
HuknERL2BvwmsFuq/NWDkA+TMMjCsptDiHSuA0nK2qW3m9XXyYqscAqeE5yJw8VpIHFPFZt/HBKP
Ei7uQBh5OisQnkQYOVGQVGsbz60FaAXGDUEmnXWxgIotx/KiF77qTkVW6Qxm74RHQWwgrD8G/1Zk
DMhPp5MYFYAzs0vNISB1IGnlYuBFyYCzs1JGaCLCUf/dtNkhfMPZnNFAZdR9yv/bpKHTB7ktzWdI
0juebdabnb4OxyT5JR+vqptRekAM95/9O8uBjvUye+arMLQJn9bBkOuUM6sFYQYkZq23DC71mTLO
kNRmgjx+fo4ktghtGnOopQfYbg4d8AIGZ5VhOiVoTBR9urluCmRmdPmGcsf/pvdTYoC+QRS0wPX8
KfSagXX4h3pV1Q2A2j6b4nwmlnDPKJzSFfSK7OMBLuj9eDK9yo2j0oBHJl6PrFLsl9vvglR16mey
fUAjbzCNYFka1kY6MwNx582x3ozyAIE0zpjqhnZH0LNuCmWWAmG6nhGPZJK630a7abMSYS0MxscW
L7Y64b/l03iPEp/d4SRViI6CjSgfC0BXKHtM1+faknjJY8Uh6fGDg8i//B27N43muPdvXPDmSAuM
uWOUimlPHSL4MnjPSkTB3l7GTMS4MU40/YIVcunyioxkZhWxIWRlQKSMjZUH8s3qfmLXjhkyJg6U
BMmp+lojVXXeNu5GL2FtGnPIV2qbv5BShcII1GkYJfYbj9IA244naoT9Y326MC7HUiJ6x/m8wLiJ
IoslOScRcgiI/jZ0Kyih7xBVy4FxjyFUeNCwD1cWwe9PlgaOpoxv35QUKkraaPn4vXaRGh+2o7We
AU203Q7fFOIBa7xh4NiQzCpk7Pd9Np0CvXSJBgotNQ0sJj/diBDYzHuz1ywE6C94V2p7Tve6rAQr
b1hYl6Z82TgBQu4GUarfLwQR0dlSIovoS4lFSToSldoQWtUwWTdhx15gH1as+VzzHAs8T6BVYWo3
+bXWM32tknUm2P0XyUzAP0lb6yJz1NtfXXFMck83zvNkJvvyf9+hgSzevapsq7tmegHaRzLoCY6X
a+dIXgB6/eX5aYkvYPAlRROu+uHgconQuMB29Zp5r9swuRueDgVgwBNR7nVhcaYZUn68G4nzN21u
E5+kIc7hkJsygP32cU/n0OIRyWXfibkAnNbkxzMsZMHOwqfOOdvdAK036n+xenPJEx0zfI4bj2U8
wSza4lUiOu/eUo2EvWuzY+0oRBlmyBp9ewq/iPJFnCOEHGfpwQB0az7MZ2RGkc+yAHpXnNszvL8X
QPD4zQeUlQKWVg3vaYg/fHNqjUwo1zutpDznl3sfNLxcvD/AmsS/C2jfDIlb+3fu7sGQXsLp2fkP
lL9JsUcyNXd6nmKF1mHQJVNjBnj/9uSnxgaWeEqnoCCzAXD48x3MBzTrN8gSa+C6XEd6L/mXIW9x
JKDEhv8ck89gUmbikaKSY09VQwnQGjvFgv461rW3d5LFP7OQh7juu8mtJCX8slhgjIwsFQuAO5Yv
lhrpat3nksHEa6RMHY5n+Z6ILeMx9RxTH1sPm1DfF70F64HXFjA2nyeUbQEBjpQBLxKgVJqcKf6p
DwFmcaGC1M8C8H1LKryc9diudforLhecf/YD57dS7RaHhMcEA4/i69ksHcn3DzMhc4wsDwvAI9hc
oi3sSrJQdp/p+yUaknEAtT6BaPk9eO/fOUUXgHnw/9EGUayktQN40rmYESpYmsdi0PbEGK1fLh0b
yKV4BVzrjcX5fw9bHS37vFazaamKMbXc1pwkGtNMGnLXFe4Oub9ns1C9xzn0e2eU21N7sB6lSKUl
MTKIl74NhK4FMdr34hUP/6UYaHms95ZszLFnQ2Fnf775P0DC72LjDn50qCLT6pNXpWcKDKpAa3WS
GjYO9Nfr2l9UNfe/X0UVsO3xJ9LG7wxv57qj6ONhwhw6/UisZ1FfqyOUfltvBFbIM0qyKIjk6xj8
bpVC8KiiRsZEzWNAInFObGWYaFpp4Bq97AKpiuDqOIImMK9UwqvW7+zh+fFbtOR3Z56tlGOoEjDk
/vzOUJugvjaJiGiGinSovRLJgORZXHy9DeFiiwRAy0ir2SohIhSFYa2/uqwINbOzonT+BR7YDZk7
hIsRRwgF/4B/qPJRwPGPU5KYwiYjSy+9gVEkDzz1pe0hWSlZyp7KgibK9+kJRpD6IpUKV4SX3GLA
S56lEPGd6Q1a07lvim4Ad3FuSJq/x6YM6nilVKO3tNjKzkPE0opOpfe+8vvMmrZfV3Zu0qZ1ec6o
XT86PpMNsE2+p7JogNSOZRhIhXYtoDV6xDOyl4rC64CMnfVnKzrzSUiTiSt+KYPqqjVnAryHJ4l3
QChuknQ153vUo3YuY/jqQWTmmFvdC9hDWfErbmWyyLKbLPG4C+h0EROtHb+St30hz8KMigyS68UC
0I8ojqL3XlkOHq2PaWKYt2Lwyl2+nP2FG7BdDIe7xGFNsNlu3O529YUwOjVxsmr4/JpbZkPIiZwW
n3lpLzx5ScTSvaq1rK7jXid4gSp8I8U3dYe8O5mvJ2f8/guhx8p9hnJeevwgVrxMWwhmK26gFPm1
ipxiqZqlOAMjK/hs7p8qW/198Z+N+DmKH6Dzu92XLQ/pqsY+Ckpy2h3MVmIxeFSH/ZB/YxofSGvF
X6TIjP5SNZyY240ok/yuG1JUSlIoeY9Hld8LrspNw475ttKp1GCDNbAh6mxgAiaCYSDbgOTeVEwl
eC6aSu9NQK1mqtY1gl4mwvGNuPBiywTHBF6XCiAC8JMQagGB1JkHPkOnE8gMSenw4zIZ/9q7w/vF
dS7FaVwRTDfES8eiliJx2Gx25TGNRhw7NCoYD+QiGszyRPoCTEToV2w/dwLVbYDJGqpfme+8c2NT
E71IP6CucRwE6pnwRSRmv431QeJLYqtnyLJbTwravtYTksHHRfsajVDO+2FO4SV+j+IrkPTMp8LY
ssBjj09HBaPCZkjqNku+rsoFuqNzZM+HRNwuROSkbCDAe2v5tuF6wAabKJ2pAEM0UxfV0OMzpJG2
4uGSQJ/kLi+Z3pBtktqXGsDHJ08WQxeE7aZ6y16+5HsHpBgWHk1M93Y76ZhQ6VRkTlgcbHXthvuB
ttdLinxqKDh2AT3xM1fv/EGHpmAhzMHHdrLh9bNF7wiMt0/k9ejhoSkODxIQHLR0B5K161H0IW7E
tr4+cZLTem+Bg/pNU1EigCn5IsrM8JIclNF7vLCT0GNXNju2IfYkaasr0frk4seoG4tkV3l22eZe
QnYW759KnyvTPO4EeNF/H36dCOHkoX0aNcwSK8Yqt6jwQ/UPKVQfVHM5CwpZ5SgzWG4edElA+qjc
GgbrD6+GFYYEPyawMlAt0aKeO22ZDZ1N0lachKBzadLM4d9hzYjf6JWyazSsYl5EG749U65Yza6M
CFHrLQNzkYonFmFv63qMEGnxe5I7n+UCfbro/B/p6aOXAFFKkP9jgPy/0pFW4EFzawiQN2e1CFmZ
0+QoGV/5OcqJpTQ/pmVtJm5viGICmxWsjOue73hKWJl6Vm1QiMA/oOqFxd6BHaxrfFd4DdRy7Qdw
eoGx8AwrOsoiEcbv1ff62nu+VqAVsI8WpDORKfCDhSi1w+ZkqyDA4kfHUbRxCVIGBQX1ryAVMrh/
OUt3ObsQR7MuL68tdyk9TO6YY6hqABfOVh/GmkKM4F5p40YYZ3dwjhprPG1UpoxfDW4Bfk3YbjOF
DzaLDs1lKOeTURJc+ItslwQOa2iYpLyTQgOR8VB11p490GSn+bxGaUueY1hEJTCQG8LOBDY5kEc7
wpD8kFF8ISmdXElrbiiPnOeUg1qnK69MRZdEClp/jks+GQCxxBsP0AwwEmv7aF+awIPrXqtKSRWb
VkYDXKw8tByNPyfq/lMtokk6jQe5S9uMg8uA6FrnFpv3+S0v7HUiFfKs61Ff7nLZYYlX/3NNrUSl
CJ7GUj2YRBReRlN2ATDv3ks0ohetB+o5n5m8BdZ78ugwhHFWUU7tynMvnnPvsmoivYGMYGZKcU6e
GkF/Q22QasHbndNrUdJ5dZ8mUz5kKEilHVx5cVt2gk+XwfYlc12pQ+oFp8EuTE/zXucZZyq/1jL0
HFF9JlhLax+RhlSQMASx+iovQkoat6b/wT8e/SItFpUuYeUVQK/GT+3He2Fcb4MP/wXGCuByiY3n
aRsVERYKeOftp91Tm7VJRJ+09ns8VnLJCSfM+zu3zdmuFqJmeg6FvhzBwOMBrKbyC3+VWiKcqq4r
FhhCq/bE8UIvaDVaUu67pDnZR9q/bquTLQoFIrEuSARHDHPY2bwUKSiTcJIigRieDr2+vm8f5Xw/
zJqorHIw0G0GeYPlHf3sCqJAnefgksKxLzVnxNrg5jOQLK1bMiqfl27pnPxYEjeDSFUKhNloURrB
tixPgsvRDQTJJjQpqhEl1BlQzSiXIcU7waQwAbkcW3XuSZNBSlxukrY52Q8HtttrUCJQ2Hp6LCms
7GyvUpYi1v9e7aPGhFnxeSAjG4F2RuE2d/oPcRa+s2RPV3FZyHfHGJJttMivP5bAvg6D9uBrbXyS
3euQdCUDqEkSjlVUNoz7ZcxiP/zcCvL/7Eccq5NgL+RXRpqqyWqII6BOV1kfowCJupSt9YKucLhA
X1tydG5Hvue0h6Zgedhgc+Oa28lLo8BcQdMYYJ7Cbqy2Gtsvzey4pdSAOtXMngPAabIR0c7mVJCJ
BwGo0Hyg7pSZt/pI7BXg6dQL7ttbcaBpfjLm400hfcyN1F5OxKZ5v3U5H8txG3Xd8RD3PIbMbR4T
FmTrQcynK3EmD6ZHVe1qGCDCRXPVAhgXsb4YpuobHhrjI2YMgNby249hz8cpW5QGOCSVeEYlSEdt
2NGO0oQ5hmOHHX0wVazuoYf5kDQxItRrfHQo7+69LFAMhHoT6gKjd+oDYxgkJ8grf1xIBmYMyqV8
bptVzvgdOggu5b6/EEB8BcvXuWY2RDtB8ROmM83vLSbpoBC5PoSTNuo+HQKn0Gwvej5wvZu84KzO
Mlru7V4t+AKsrLfqs2nGXjJIMQHZSmLBmpkBzN54bg/+CIrJiOvoZ3JE00HMjGi2SPP72oJ5JmvM
j0TrtZe5P1QpZKgbeElHkiWH3QDp/4iu7JZz8Y1CN5oPxZjM+E9gPseHbmCshdzXmaPECoXOQQ52
BGbf8Yn2ejCvWGmo40XV6l9ov2dTBZErR12Cb8z9zs0IjyVg6Izw6rDyRRI79XFxTGHScxW7jJdN
50cFziSkBP51TrVBdFYrwXlsLHpV3khItoM7D7pdL2jEDjGdEfF9jYw9ZlwOsx5hRzDMS6Gv11pf
K4iS5QhG8D5gEfr1taja5/XY1i1yBMha8zGB9QxyGowzTJ1zywkIt8l4KXgGibm/7VfLFF1RB30U
hqv/OsmxH9NRvDSfHxoRCIRlhMXMw1u0A2lPM3Qtp85kvM/3nTZcGxqPYfaLRomha/kB4rhkt+Sj
KPVZGYJ50GDqbHgbt/FJo1MP2k+sBdC1DUJ/tPf+DPQlYKBYhwaQj0TzYwW2wU08tLCiT370rG0z
aGyE1ZPlqbhRmFPiZ3bc9DMEC5qTHsNp3v+lMTgAc+w7Ajk7GUo+qJEmiiivqlNtOYsjKaod48Xd
SI5IbjEvYH4ToJYyDhQiEF50EcoOJncdDo8P4TF+mgDoBFomNd/x7ACduf2XVfgkNqN6690PSTEq
q+DXvXd0osVVBa6KGvgYlLHDY5GT+cLjv5O6mqWa7LcqQxc54NddpoBvlSV952qhKqn2/Yxjn0l1
i11GT414JZvl2vUj8WIjFXaBItUis1tZQpgXWq9uslpcTAm78VQ/PpI9X4xlcXDcSKFh8IPvtt66
OctJAssFEAbY1N4KpjCRGQoGc7di6jdgvBnQ1ZYdBFSeAB19tqXwOHII7qjL9LiHDK+DyouiZhQ8
WjSxgWGOXv8noEZy5CFBMb5adQFr4wG0UxqYficfSgVLumqCHE6zZOmR2v2ceSaEVgZZAvXVnf4l
6EWEgLYDT+5FICSwryU6hL96gkkns0V+jZak/jzH+SAhOgS1AbJRVCYKp9ThbRCbOgd8V5AYhRE1
Q58DwGlwSWrV1OZkt8xrhTEBYkGtPOikwHULzPr0ffpMNAsECTBpeF/NPj0iss6KICK4Q/KB005e
Sco1sIF5XPa2jMjpQ/7u5ms+0cLqQivl2HoB1JURUrBolv+56+6hnO7RFMvDDpsHU3+DcWNl+rE7
fON2bxBhrdnzw4kfqSb/+Qp80DsErhccRV2LWo2zY/pjowEasIBImkrx61eKefk6xcPAbAzVFB25
YjdYUPRU9rJ5/BQ/zGXx60Fw9kR4KuFkhmk7bIkz5KDOkFx52CM6703PwWZxQT/eoU2xDIg+oVTE
485s7UBWczeFX2AREvfJunvAkVhrBTPpJsbvqgAkaJAo/YIy3+WFjYDipQfPBmLJeTOv94u3A0hh
clq/0k1aFlLUojsLCeTw9UMFEKBP6YgwNcla+EHYeycPm/g+ONgt/8hma+2aGaVsaaD1Oo/bC9aT
FaVCUKRkStpg5/yrxBOQT8i0ULrk9HEq8mJ1bwY7ZLL3aE4/BQWKoUX/ugxRgj7xubM5zEocQV8y
YtUrhpe6PzwFJDnftWMgFVMbVg3SDmsruPf+P5X1/bsY0k0edUsx/qkmCQAjTsQ56yucJ4rIGFt4
lJKbYipaZv4k05uy8m3trp4iTHwTFeOjpESyB/FVNaJKJ7f4b79CnTmtS9kapkAAUCN3QhjymCGq
HPYju/x6afCUUFn1SkGO/SyIP5/HMpGHb5Q04n92EMaIZYktb6X6mLoji7E9T4rklQhR44dI7mkE
BKl7Tdd0YsLZKlLdh2uaRxsLlZR16l9pyr8D+zEgKlGYFiuaQIjG4YddjF5XzjNXHo5hv+HqrbTn
cUAIBH1cRfozadsn8rYCUUmpyxOqmYu0kaMSPMarFf4HDKRDDR1nKawGsAhbNFHWCRhZL2J1q87R
xw2KgGn3d7W2BlGx1w1k0TGlF0BRQhzrdtugR+Hm+zJ3V/wiJvpXkr0/y22u9uTkpHTSIQh+1aFp
MeTCSLLO/txY/pdNYtcLG012FGDG9JKs6WJEKOAi80xRoD9z1j7mEKVwrOmaT/vyhaHKKdzk4MeT
S2BHWLxUGFA47b+5Yzsc4UkcRB4UEmjPJ0BwRdxcysXgTz+mBjqK7eCRHuPHPF8H9vszJy9bs3ca
nhPl41/CyZBF1hNLOwAO6jBd+9HU+H9GBgxjJZ5y3brLNsfJ+07jzE72d2a03uH58SaNO1wQi19o
xwmXhxgiKmjJ+dorb7h1+v1WI0E4w1+7pHWbWeC4uOhVwj51szcvUH/nApDZzc6jmbtn45TQnbC8
m8oSMmusJ0ISv76nDmspNrYK3bSg+OFo5D/IxoYUieP3z68KKHdedoej1K5D2TpTLnR6pBnz5p2F
fVxOmAtTxu1WeQbfheTKky1lbf/j5bt7FH8ZGgGYYDKGCEqHOWVDGPMzRWRX5wm17z3r3Amtr7rl
lMdZZbq8JfF1fTnqiCy1PnBqEQqN39PXJDtgRV5AJvEuVPLBXjU6ljQW4w8RWV2K55+6qCukSPui
uQeoUwZvSh6Ary/sMg+v2w8r6+ubuSyo5jq/gaHwGNGW/L5RBSssoDi3cFesUM0T6zvYUrkwVcwi
5NbfBWkajw7iydzjKQddS+e1J++0Xzy8p/1JpokGkMsWDVHfXYjFdH/BY8LGef2/Nrkros+BEaKb
274G0a765r6esqe90TfFbe13H83n3E8C+8WYa7ABMiR8gBPagT/QVAPj2ZSEQmuz8KtdLHxLp+hz
tqoL5/l2AYZfgGJbEnnFX2tUHL3i8vDyTJ9CaUDlm1NraKz5tokOlTcy27BRX8hNrLnAjDWPlUk5
jsz2a6NOtOA7OYy8xSJaTLNG2BhwcRxy1hP/OiKuxPqGSzv91ahoeEFZBP2c6XvSYdpZL1A8P7av
rnniTS/94sF80rJ1JaSm4LdU1XVzqvrNrb2luEeOBGYuASmTpaQqE8Yfaj/vVsgZNZMPG4Zmp+HB
NpNX3Mz6nKhEX0jdRk2WYTdYQ3Lu9xaolJdlzyeeXo1dmlHPxWOvMyllXL7CK1L21kx7SHmUMBca
qoiMxJgOAyLSElkAuHEWNw0QmrpEtdubZg7GC/QKZ1p6FPZHsNbgN0lZU29P6Hj3tS6ISiNvAyzO
7336Q6szSemWG74MqlWVgxJeVk9P07ffCFffFJPYEU9poDpc4lpP7tYD8M4f0Ox0M5OFBWe31SxX
2n5ITpolpkZrfTXAdXwSYYTbXHrhbrUl5f3mxqx6iIvJIU/EaJ5iE057t3o6JwnuaHITbJVTKVjO
rWlyQkALgU9vUvqkwZ6jMMSMV2nitB0oqS7GZQop/5Aj5dJXor+CNK63IjKfVd/jJweWkDevh3n9
rpA/1dWjm/67wgXuLk9tK30KqpOmakfptGVEj0tMB+i+0FCmpLVBLqKpmJFeAYzSta2ln3kepeDF
Nt/fn3kAfDcbcnN6nqllbiadS4IMvSLD3COW6OMWLi4Lr2PQjl5FlwPp5XP4cczmb/VK9F+aAlxp
e5OAvDeIdRu3fJKpZELuMh7fdBBmqhVHD4+KZOBX4qJ4ix4as4Vmn2cMyMOkw6mSqwQol50P1o+p
R70JfOQjG+UW1GT5zJPOgAm8iBtRbfwU359lagM3ey4KGiDnB9/OLmgHCU9ovVftON/uEMNPBkHk
zAaf4paPX1hISqksWU3nEcUKSFuFhjB/LjZJumshkCmefmbwgCC7kSt4Sud+/v7PCeIExmxW0vEO
fYU4hPG1L2StKyqzmDpeSOh1RtbO8PeAstJXV6jrJcU4jFbFaK9fRnfaqjbbSP/H3uAakEfzbwyH
s8irEcrQWVhFzCBLFnhd3A5oOkvn3gABJktA1XStXBy+4Z8BmzQIZTr4KOS15eYPuaAfKiKxd19R
qKsUQ0CMGA63+YUz2x/OvjxCnComIxeTT4hwuXF9o05gkAQcTaCyY/xelAI8+wUrGHDpvT5iktMi
tg0dU59vTJ+lanOhw150vOoxOeOvp1Rb1WU0SPlJ8D13Bd1t+MTL5m0FJWaelNNZc4f9sYuiy0rO
Uo93H4hHdR1EB76vfYeWT8lVCztFxcO7imtxDv4c5TpvGNJmYMe76qGT7FvYCP/uQkFdubNQ2bLK
hOTCXBs3E/sJ9qMijPQEh/xhNZL3P1OgC7d4NZQhq5SBDiG/2j+q8lOMOEB942WjMXAwnmFwvztW
pCvsiM1vcP/myeJffU+2XIbxwttbWg+NEujyP7URXrr7XoGxzXiCA7puXQqJ+VKjyhplzynxRDMp
f2Bh6cmaK/u4hGTVcmsqPdmzWZv/GpDdG1jqCh9KzG/nAHLY91Etsb3DCvv+5qw1BGGloYLXLk5G
KeW8dVjJUHlj7m4TvaeaRyR/pgdqMKyQDJD77R/E4f404z5H0WfgxshEwXttsRvkKw+Qt6PnOYp/
mK5ak8mmxMjtx1YkdFdbRy7XQ+wwPXZCeqR4PgfA0ZTLwoFrTSTiHAHrclOf0ckZrejlz5TEpf/u
wUOLSUVvmy+IMoMiyEi8yDh0CWPx6/9s3Z0cc6a7VCn8bldoualzQ4BC2elmcZS3Cd4yiMvLBkhF
5/muhFnjXQtezMmgJwCTb62AG9l//GlDHKPTPcW3JN71uYKbK4kGr38UH+laRC7rFyBm3XAFy5Nq
Y4f+a5Uo2pm7by7QgauyCKaOqtWzhcF+BfC3GHFaV4UnYjzu87rAxc5apXzbRTrT6rcgXiRbKGqP
3um0AAnyTykcFtQuw9FPyF2RWD03JjMQhNGb4ai4LxiyseipF/23ZuUr4ip8Nz+VL3QvpoSiiKog
HdZktCA1QjtgFFPB1Rgo03Xbnxc72pegAIGfPnucHyDVClWjScAvfYSWaIhGqY3KN28lRKm8qgV8
Ye1vHeJKcjnIl1V+UOpeepdgchJt1525dhoobdtOCrrUj9s/h8G3/GvoLDF4Lp70Dt3k90ei76sO
/2sbWI3n7fbL1vLWkJJk657emy+xkpIyOcm9LBqZbwSzSzAzH8MUGXUaOfJ2s2P/SmpN1eVzFLJy
dn5PR2BmJFTRvtWcq6ftALN8u2X622ILUSl0dG0FyXTncvBf4czS4VaPeohBj67FgvmSAb+Lp37F
eqnVz5xRSS0BupXf+tLwYlHEaEWtp1/f3dRaJkS+Tr/Cl9W8x4GHot0+sd7MxSaSjDpTwXTfB7AX
nlQNHlVj5OddB17/kyY3ptLOLNtfdiiaO9mbvoXJYpWP+t9k4/hfYND0Rka+hKdfIqVM/lAtmbCY
QMTbv3p1cjggw58QFpCL1qkf6cYBVlK5IYNNxde8PvTIAEqJyeDoWfc8vexyho9Q+2Mlibd7OFrZ
R2LWGENozp4tux8zH/D7J+F4cPAxqZes922SX958k228yWUTdTGX0nJsHUcoeTbR1hDQHEWEH6Tp
gY4Qa7BNTmSf/5LrRWDGBzWvP/cCz2rIk99dvKUzHqBW9vHU+5uozX+aKEBbIUcwr4QzFewglaoH
cWhMNQb9S/E3gooywd9a+BY74DeZOkGovRU1M8USPcgSf4U235ap+66kkdKN/MMPEtj/rrvYunJK
vZtYmC4dKZah11D1vMC1+E8fSA5Q5877MnJftYvKu/sHcMZEGpW3x/G5MaX2kIvGyb/RxWFfkcmC
QEnACG2+83dnahlEvf+IweRNC+RtLhsTN/t3CDuEBBM8Wkz8z6Qh98QWix6caH7Uu9MzTi0HJJYM
D/xGK5PGwka1GK89R2AzByUOwqTwwvzrN484zEH9GDbeFc0s14W5x/4rsajTJb73Js9DFsQYfFEi
8dclKwuMxleJImxH3p4joUcmwH2AP2T2tjg6NmdcEwyBPm8iZG+tiej0Oaw/6+nGQogL27EPozuj
MkTxjGALE8nm7uUSCFU6A0C6iWsDTlXJpmHk8WbB0TEJVOa7c5Ncm/fp5UQhz/LV/6M08WICPX8j
WCGD0akQrA580/mI/SBeNiwAowi0EtU8MNlROiq0Xs1e7LC5IwNbBDB6l/ju7ENxoAHhnDhl7uXt
os/BVWUVyr/8R7+AInOcEwtWgB3Qo0vzoNmW2FNxClWcafaPP1QTf4aorytqtrCCICVoBPND/vs5
OJyYRwwffDftG3SbZRX+QE8ytdzWn0d3QaRThb7rHGpxNeg92+PJyW0nXbUwds4L46Ot3NV4gw2O
RrW+xgms8x0vyglvUmSBbtu9P+/7XzmEA4VQ2aYezniCQt9IXxWiw4KBjW6Gjec+JsppE4+rmRuq
sEwT31VhwAR26YIRVTcNB3sIx1+ok9F2FBY3E3IFhzZ8pmaREAqTjcPReFJANkscF/OeP613hoT/
x9xWNnNqs7eOxgiTJ6/nCL9Bb9iUN0j21nzmDsTszqmxLvWVwIqXCE31mdJK69XaCBTlQ7+zsQm9
JyoVvobjiK5nIPEO7E9CmNbVNHfbbtNnZXB+orRDYaOfgDdWIAKPw3ceXd6DrAdFakozTKKYdstA
zZF0eZhBYqWa0UF8G6zgCZLbJe6PMeN2fMO+TcC+ISNbYhlpjdynIOWQ+oeav02nJZTjwYa2+QMo
yJ6OLBmy/w2LTfCW8AgZy3602/9jdzGvBjH3ng4Tb/C/7rh8c5rgyrUn9K36UE94BQAGzxByyhtK
zT+9IUUNskSKVP3DXC+YUKeWj1hcI8HGl5bq5E4gq5kRYum83bp2BffZKg9CngvfVFnOKmCzSgHB
B5FX67UhdeO12yw3uSV4PysyXgfhrfSWdnsbpNLFwyOodjgSjmi5/wYKgy7aRcgi9bTuP8DZLmWY
+0rUVdR6JIPwqGK7DUc0vdRt0fjzu9kq7dNs2hhIKH0M8XkHR0VtBJs+Zf/MqTSfkFM3TKjguwtL
Ufsy7a1DPAa2Kr98mFvslZGD8N0RSNaGC0+88x0OYpHkJcAWVdIIrwZth2Y4tQRN5v8JH6aCdzfQ
fCjfhH9QV03Sat+kes1z8vkuhZeNpKQaH3lVSg4t8dLFTPmQZARBulZmU21sAOxPsrCG0Kzkrp45
e7ZsqshhcAGjD34RTPpdwUhCshq7kf5zlTvHGPXIxxOqATV6N2GByr27hPMm3CP8KNlMSQuCZN9g
A2PTdmQNDy44NGBHZc032w5Ge7QN2MPx+W/omKnSSN/qxVLTljJOOSchRswutRzQVDMgWVHr84tw
lSKDsPkNAvhgtYKyJnkPNhnvGZEwCUS6FK+xM3hUFyeh7KYY8RieRgXOC9apuC+codh2uZ+6B53R
P3amCOG131WkXFbgAYAM7l10NvHI96wsKekVVgTRFvPF9wzPPCgj0QgCBeivcnrFWeV7SvGBfVmU
+v+IZJrfEgF8/QRj7rEuW+hMJ8/ykQVx72SIo5SP5OeQ2OJCxCZCRb6py+las6yj1aofyRteeq0B
23bolrqFEns9KatuuA/OO1RouK8uGTF7fZn2re0qPeqJrZDO2GxJxVt3A9CrVYP96PRo7g4n2Ugp
JUDLuLcvMU/dizTQoEljlEBhi8uHLxae3K8hNm4GgkrQqVhBwjzZH6mzvC81f6q72R8Kv1RETXbD
hGZgX5Mpvr3/RrnWxXrSMEiN1YnP3Vw6rxL0TAjGZ1n5yo8s2PhLlpXxqBAFClfWFuPP9yz3bSHJ
/bueOEyFWN0IimxKf2YDQrrEWkSzXZ+jkRPm6soMobuXNv0UabRhtVOs4F3H8ocKm/Csp/w+ZNWW
HLUFwvF8s6WCFjMv38ni0nB0C/IlRXJBpfuUrmEM0PZYP6AZUgS80v0zxY9o0UhQKrrxRO+FnZjO
D7NOHUnMH1wdhSKdiODNiNN3RyC1hlYw2apb9OWp9+8/T03od5ph7TrQT5Xlzuv3B8jJ7OGSqhO6
hizyPu974gjA4ltPoSFW62JJ9qpAWtIN+j0jb0EwYJivBpVtileGTvqQauqmLvjAUA3d3Qed2T4N
V9tXR1IrbFldVjZAtQLxCJwwmT0wYatOrp5+oExr6oVljJXU+H3C1g/XQ3b+lrBmGKdXqtvHXZMP
9MINQTCD1arm0Ip34XEYGM+QTgnrH5gmiNBveJW/RqmZS6XDYyQ8hz35XJbD4cMDEdad5Yvgh4Zd
0keooSbDSZdasPnhuFYLh5rP6JmUH18rF2CFw1uiYjd8zQgrpiTOAV4BKNoUj4hV12jdzOIJAMcI
AaGwzp1ZZZd4SjN3JZ9LR0pG0W6t0JCOGHHfDAbegCEcUw8t2iw6vqiVQUlxAA1jKaXTM8+BcfHD
zHTAfZs0npmyyF+e55kVk2W0koecKqsNwlWbjINTee1/zhP17q78FoHWL+YgnPTYvpL1vr29IJmo
bvBuxnmI6SwSzg2SFZfx52iiohFUfOcF8XoLzIZC1ccJJK5cBKmWIHaQ4RRL66P9WngUz8qrcoPn
FFuJub2Ezlbu7tw8hsCTfNjNZq2MqSLHLpY7OUglKCLa8otmIqwctS7Ho+ykpHhYCz5qP9Xi3PDe
4iLjeeXRY3CPKufyrX6JxtsKepEV1MYMfgo6kYDxQYov6X+qIbkIX/ROFkKfjoNZL9XUz+ognFSY
TQNDhWoFNS4j/zihAyIBsSjF6C7EPtlo+U5th7zVrKM7A2uXctOEFQ6iLVSiuwUnhGNH/VdBRXpl
wreSeeX1DRBCsMQCJXlJ6su5zag3F9gmLb/ZIzr3A8HREy6OmlBqyaHeEswSoc/hCdwzSKu4MAoA
4k+bkpsakMe18Lwuoxt5lc5MYRw51g3I/fFwnVCRjHZ4VRkToA3rg/O53Blbh+iiDzNdpXJleDyE
SrQ8F1WTSaLQ3MLmD/M537cWo0BIoVn78OQmSjBdeHteY+qUBphTlrp2JcV8EvcDVDJHSnE5Ic6x
SUu0hMvvocGgUkVjbL/7tBU0nL5lDN86KxNq+1SOrxGjShwPCPdIk+3kwVsug7i0/3ENEUYsdAnQ
bnWdG/6qU4BXftKg2+U/l4absLyHpeJlzRxB03HHkRegPWprN7QgzkUnl2ucGNu+i/D3ZtPT5nZD
uGUiAWakHGcljLcglzNjujx5AhMgEjOxwrqfOmfODQgldGuX7NUC8QZl1sQYSvwL/NL/Oqsl4GjP
09XHFXYeWn/Wp0VrStdsj92qOlSAw1MXbIYrubdjrLQQbIBCS9yFbRSNi52a8kjvJ9/x8ohMNhhh
Xny3F83WUiD5wlDQfqaCM6Q4vtZn+ndYJOmuv2wJcI3OrDME1IX+0tQZa5hk4P2JbW5QoX3ZpJNH
TuewXWOP936LQKrY5AncZTBKTSEIUbTrFmOkOvoxf4ZN3MN7TkErPH3gYXIeRBXkrSYB8Y8doAc9
4g51jkG+fNpQn9U75Qe39i+WCFiCNhlLLlHhBOqk8lTHxgrf8yWYBgsFqKWZnz5T1XsMdxiW13F/
YCz/7sCnK9vDUlVdEEEPqgWTtLpyeVYovvPp7coNSn8AYQomXjE8vDEHI1+BS9alRb03NtgisrBx
4TMqqfbVyRx+lqWbht9fOsK0MKRh5z2Tk/jQC76MGxYo7aayPQSe+8KrnszGLT6Rf0gBv2cay4iy
sREKIoK5YuoMxC8fAdt0edJ4yG1CZD3aV7/Vnge8TWCwDKwSIIBWyKf9m0YzSRu45+MvQIMf+Pod
rOhng80nqN+MbeQM8RefYgUFVHtzm2yLgvEsCP5Uk82OeHEElgzwjvi/tFJflvzQeFmCOKKF67Sb
PWohHZIGTKEKi1v8KTcZ8WPwEYK4UJjj96alRZM21oOCK7jkhss6mrIKG+xy0w2JQ9F6cqJ7lVF0
claGP4vLvOBFtRYTg5eOHXvBZ9tZx9yHh8kizDcy4MMW5/ZhMx/84x0u0WLCTFobN+LeoeNGJTt1
PduYEqaVQTzIsbLt5FRW8K4kt9jGPmNbPqruOVhjiKStsVyZf72bBnokQhVuSrE0cHPWqCnFLbN0
TxW0D4qr2Nfc+OQo+23YnPUEUGTROBySgoCrc2W57MnqOqeAS0okI2BsHGPZWMykWrJ4aV/C3csa
jIqX+z/tQOhwFLpouM7FWGAfuf5M7YLf4T6YhAiY/UmMxmZOBQwTHRZ2tXk1AgOrvnUEKNug4l+g
KxwnctD2nrKQXUq+PML7AdbfzTjs91GAHlnHxzlTC6TjVKwIWXlBUU7FFFe7y5pL8JT106kc/5vO
IovHwb4g5zICY+qGKDWXm5+B9HDxuFZVKac6rEzGOzXVvJvhFoOlJWgnLWbpfCcPikzPdgwYX9Oz
98HKuRp+bpY8oHXxwRKZOn4eUzcve5ANjH8Xc298kFFEcV3dtnOFtYFFBqIG+xMmDx86CdhGhvzy
FT1NI24WggzaTwpekQc6314cjlShS7WtKkfNopKJ1erE5MRruoVwxbcGVvjR/s7c3eh97h23mgVM
s9ZmfybZTqLeS8veRcuV2OB+oNiZ2LzXrwNMsr3ZeGMOha3oYlFJ8eY4B+M8R+v9bNhQWjXbxRIV
3grMObvx3J5IGQkc3TNWaMyz5yNZVz7Y1hM93andDwpAuF/5uqmc1N805SZucBYR79BKeIjM/34I
jyY/zPvolZo7csn+Wozb4gyqzpcKOL5mH8kfYhUIwtuExoUFwKtidbY7zUBD51JbYX+wuqy15CkR
/IABFN+JBFlBo3bd7hVs22QAvXHjnWNj9PsFsxRZYXxV7liVdA2m1qj2vuwNK+/VUMFZGo27CK34
d7CotyameVlxsTv1kr7d6/95x/oJDDc+0ETvadajote2hPygLp02XiBw3Zn/v7IJpQuO1NnlTsuQ
m6OWcWciya37o4IC06kOqsYrXhdxg+Iqs+ZgRAqp0vpOZFPYaCLEOEkZ4IuSrhLHFWpmcngE3Ep8
QcalEWvvQwA40D/5Zef+m+PDd4/JcJQxyYX6XG+mm1PGp2Ej4S4FaoofVYbzhm3bBIJlh5OCOGgf
v97lTzRz1XVJESA7SdEglEY/vMv/f7TnQz0aPlP150cwFAueAaAP/qFLKmxznvngXxUD9gyRElI5
7QnPUZxwt+HWGgq97tcQ2KUtU/LhYfk5OlvDFMtRMlypHKEDoZXZ52ibwNUbv963l2E/p4LYH1oG
bZlqpmTi3ObGPU5fimrnZB8EfEEPAl5UXe7K15XM0GQIKoBXtZSaHjsq/iwLxj8beU6xHK7wl7ED
omsEXyokB/XBAykqVnipfRmz8Etd3fkDU8qw+eeqsdwoUDioSVFSFZcMPALSXs+IJy8OUHwA0pGt
/EE2MBRJwytkPmSg3SuALFW5L3GgPPApGQYMS4KoYIo4CbkiEFIlrGVp1Ryvs7xYghWrJlPcGghw
fmPeEb1gByxuBOoRcPQj+GkTc2GuW9dTsL8Kv7/QltfanZ6I4d8TwixQUgl+6dpfT1WTbjhDCPtx
MHQCOwJpwHWSRLNC+8EjigKbfwmuVJzO/3WbZPZFCCdWgdN8x4GQMUBghlHD3ohyxIg7LtVTI/yY
mYecerMUXwZnWOSNEnKjnR20f34/Xb/ELaKVhNKwNgmkhrnvYvoOxLcqDNjZGBbaxTDJdQ8fURR2
mFZYceFAZgBaIFu6Qm+6RVvm5GLf5hxVgl97SlJV2mr4bjxMomkYy8qnKa7R2fgp81nIjGpLf5qE
H/FCsdu10/W5EYmtTVCi6xlUX5Iq83slfClmjWHRGERC8gcR6lUvNE7DDzrGzNynkekfvEqYSQSv
EtUhf0JpZ6+/CeR8KEEzHibQFMFOtYDFU/gbhltXFJlOqyl7pBgqjAv+TCSh5nrct6FWnN5wDGfQ
5Vg9eYF0PrmGWzEtzrsHi/c3PrVHaYyPS7On+qvdvw1ERNQvwcdIBARm4xfq/KhyaTjeiTbqGRHF
SoFOMyUcFDVB3zG8dhtcznTNgVcjosPfja8cmDqo33ZaM8eTNDYrn3qy++XgFqY68Q3A4Julesd5
+3d9/XyRkO5iAWkwUMZOEhKrG5+z3t2LednuzLDYNIova+Ed8ZbLyU4yppA3hg2JnkvGbDhsF7Nq
v3EYq/QYhN25rACM8/MvCzB06puDL0PRaSLhlA5OjBUUuud98wiMmZlpnND5pQUSX5zTZkMcPMyW
+bj0HFCoFyPm4fBEaMFkcwgugDsv8MNGIJI+UZ6VXCwnArEx2h5wRAX6xQ/I2tf6OZjX9AN6RqRM
wNXLA1gWvEEGYREHAFohkXMX+vU0CMn2+2m2wWyf5ZFO2oWoPBx1zTBWA46mmVVpJiOeMT39vNg6
tv25H+Md5CCC+zXlVPrg1AagIZxXY2CIjGLgbFDbqlmKta/IRwsIqQux4HC2t2FGxZCePJwxddTw
wslE3nHlyNunELYecoFBTCbn0QQh0+/N+p4/WVtQin9ameIIE4hXkwTKDhEzfTEkuwaSbrXA6+qR
0wYtClWPJ6Zn/qxwNmsgqaJ4daS/L4DFRpDKYX8BTxC4rhbdHQFo7TjpCMIQ1ObrGn7gJDGRfa9O
9CMjUNab6mRkMdJyiKmitWzP/7w0N/fYtShkMDYjGXhp57SeyJJg3i2OdC/30UPDTMeNQw48We9k
1q3YPVVn6msjJrBrM4YSfByDDNHj+eh/7AxERjyBCQKZXsT6AHsMLZBLFLSDz6ltU+2D220cplOJ
qWJLKHkZ8PRkXHnU+DeRs8R7Gb6V2sUNEA0b7vUrAzT/OKs/2sOEqvIjoBEA4AtrlW6v1zNpI4g8
iV4WwKu6o46GwNy/RpNPLzmUU49VxZ/6zBefly717Toa4ajd2LgSNzkeYp916ytDL9YX7iB5ex+z
0edN7lVqcWB/aKcOOCpEoY7KZVNWMipTr0R9N/FQUyVwUbJ7OsrTQBgeK0IgwcODY30+tGahphFG
Pvc4PLbSE5tVu0dLtJD70zRuN8UU+vRsOFGa6thfmdmEP1o4SJkE68QJ57aZT+x5DtyCmMXSWHsA
FrUhYzM2L36IJApM9gxv+l+GjNFKiAh9DJcjeduq5WxKT+XCkF4u8uuSWLQzPQIuRnkI7P+WTbbQ
5U7WEehfK9//cxwqF0DpQeiZuSIRXsPHRmzRr29xZ2k5oXfMoehzZ+7nBWhC85NQkAg0xXpTOBa5
Q1J+MO7MQAUE3+EOtRIo13JPphZpRJGh6nOsNbG5YvrdizJ3Nb/BlTJzbZVa8AHVk2pZGj7mHIAi
/1l4NotCI1RA3uJJA1WHShZ+A5/JT5gn2jMwB43F4g6tT5MYpCGSwuGXd0p7rY6A3MHSQcvFLoEV
b33kN7kJtFUDxdVgaq98yH7bSQVUNWatVexJPZFAefsH56qf0VdiJaTN+nxRJQI5qB3lTBjvosZA
kpEddfTNbvNC9fkIYYQQz+WCFTQZEFsYWy77EPa3JEmVRaby4v/9xH6ZKJdOZioA1aJQ/bCZ/XRR
Wm3j6r1NfJZctSTY02GVkK7uV2FbuZgk9zxREOSv889qybYNN+DgLl9H96Y816ymnNuWnPXAYWsu
QowiGuohK12HNytDb6OeSUCV1R53gzNlTFbERG0dhB4xhpuh848xkcJxPGzckb/S3WlWEfTN6/FS
7vfMaXAojWzfCbinQ6J2qR5ks9IVAtSC231HkPnFzTVxBafw1SR4lgymby75imasp3dZwClT7Hlf
q1uufgwxzChCjS3d1nnAVSoFOEbvUuG09OFYNmeqybOLEnqG+ciSdtUQ7nDvIKEoOZijLjlJuf5C
vAR05ebpwAuldZ3Zuf4VAWAqYUjxqktY4l7ctfpAz4OuJxBsg62XKICuAJWaDOpxCJegjCV5N8JH
Th3H/4ODedNNABN8xlu4Ty5ulODrJTO41cTv5nZEP6OW3xc5FDpqrML7CiWeEnO3kWchqSilKlyM
bjK2eEXA77EzvcFbb2xqfGtxD82P0Z1kqrHBnlESDHU6JXgiOGTGNHT4NruxrVf63O0CkI/E2RYP
MIzaPMx3zKuvx+W0F3HSrHYHyLVDWoTvxMlSeB9nP+taroGtorWww1bArpX398qFBH3DAwULYt2X
wJN77U/dOrnO/CRGBL6/oWVurzmXUs4o4Juthrx7oo/8BoX2FNO4kffTsROsTlYhy7NSMU8Q3QAx
aW49+kbDR12mCFCo/kYZ8qU2k6oQoj26x+sWcQBPA/TvO7fcq9QsQUiXXZqiLgJKN/vCOPuM0Wsc
3MZYNZ95LClpx4Yw0072okhzc/kEGDnvMxBWLNxTq+4UaSrMnyEQUs7uak6dSawdHwMfyX6+jJVQ
wW75ScH4vtrco6wOWfNiz9cTtxQP5qzE0NG0sCgXKfk+vc0MA/Zu5Bw5s+nmjynvsu26n7J4oTJU
zn+Vd9pj2dKfTzTJ8NtcUjIuYRq6ru+HKSkiaS7Rt6fVEZ8mFIs5wQPfkBJ0knj6HaqnqnZXCxtr
SbCzf8GJ5khrnLvkLh7jfJBaCLuTTz6GCtW5Epm9mgzszgzxQj4zjVgPBHgHb9S9r/ZQPIaWMPy1
Q6TgstycWayVPrO0MrlDXnqVUaQPqgjQtAkX/oZLut0NMktNDdaGraTFqFObtdaGVpYCPCN8gHSV
BxomltXHBWpMFgpt/WjsPT4Jqspx/tRQ7+dPJJAPYSNw6dkoVzPWqZ4ZYv7SaZF/fVxb7cKxFj7p
9gF8r1JbUdzKko3j/1xwm219Sp0ePum73vCqaNR0F7yEh2mUeOXSXwkWQtlOd1fr3aP/2mTl/6sM
ZjIV0uDPylbB4aTooDHR0qxVGtAGIX+dX0jJ+Rmy5noN5zfwGz/eKN8QC6bZtvaSwdmlU4ww2hJZ
dL4hvoaACwY5i2zLt4OuVpFHqz0QznQbjZHTKc5lldsrl/x01VoBB30iABolol1wUH49dXD/A8/4
qC6v1fF+t+VtoHDCk1LG4obnj7UZpY4t8Da2rLBcvHnWCAwWWqNi7mlQV0gREFYtxv78RMxDxW94
vP4LnW0Mb0Dmf84B09Jy0B+qg5svcbtwA3j10t9Jnhku/lY2UwZO3BZh/rpSQY1RUyDCC+gVzDN+
eQYGiuRu3J9dm28KtLk3CIZSOFGu2k0fsPAvIlPoRUj5xzayJ8kHjPXFklhYfY+KqPSjeRffnfr9
H4ckmduCrhhE5z2h5Mt/mic5AxXzbEP2vQwslE8GWOYjzUyA3Qo+OQbTUeHok1MmwFTRGgEwpy2g
X5Bny/Sr+398yNFzWnV7cfNVQGOzd5Zw9sFItRKNexAE8nyb1/l2BQlV01WtBhaxPrxS696kAMjU
9Ku0FURlYGtsL7M8Lr/F+bfjhSYvhvx9sNeHjMiD1y0ZAnczLa6Ec5ZhnTsQ7TbJudIKn7ofq0fc
zImUkqofHb3O/+R6dRcJhYs1O/ryV9rXr9suOE+TWt1Lnyl2sUhXjAx0pK7UOsY1mGOlY5qIfG7z
Q+i6A40sWu0Be99k4xe59JirpY5VAv3bubCREsweTWJAZDJJ6ld009zLKCZq9n+4nOjbVnhiXEy3
Zw+RVWnCztH+kwzntxsdAgDgZ5ghNA4paG2wonNcw3fzMZTdL/d2FUZFq/chpHEU9wOtKRopxgjm
8jhlTl2GPZZQpoCsazvnHk+lWyLkfgbRdsziElnXKbxODgbmzrrIvX+lDI55XyPGRXU0Tzzg1rNz
92rjfVNyQN83T2bt9Mh6PZYX4dYuTrPkrm7Zdiunv4+zCEStVVPYm+oCNmiMbZ1gVz4pO9FC9pQQ
zghOdDmINizF4FL625acjpEmyHi9cD1LPJ+kF3Cak4lP2tiFEb0p763zwLdMKNMCtgV4hdq1kH93
TeJpS1BJPsBfHK2BCm+cx3dYdAeDPNTTtLePUbMIkUpiXNJ8BrEPqDhA4OQAv/LJgiGnPEAU2FSf
c4b+J4gpVgOLqTgoD9AgPKlGzE2kGjunjt+iPDzCEraz2Q39ox+lwcDBqtKUjvbrv3LzE2buq9tS
t0x8afo6A2pJM9jJKZkjjkKaiIN2x4nU/oZrU33fcpzC/GA/Lkh/SA52zGEuWl0unWFq3aimGKYB
BqX2OTu35wkyOqccYL/Yg6sWQvFaiUb4G53+WQlty2ypIC8l4RIzE78E+zIPHzqsFRT6wfrBuY78
69yRYmmzOzGvyLtqSVgFmBy8voSTVfMm3vdEoYRU3o0TVLHYEPq+PnjWAAe5D9/OgkEMEuwWuAD7
lGO2ZQ6TPJW+B/o4WozOh48XyMMrzXcSCifU3mghbOvvSNqzJH8j1sipI4E2aOJug31MPnpA1gdt
e4e9ng0U0OME1ZLF+UU7dn4If0oA+WZdIFDK+gr2jJv56G+A5Z5k8T80d1LxYc91pv/6sDy7ek3p
omhyUyUAXFiSLVzhGSyX6NhWWWRKTGvnIeTQcyEOCzYtiStZCPjYqtJJS2w9l9jGuTlpfd5j1ELk
FhIiOaAeF95vrxS0ukHUix5O3MLOhSZMkae5uG2TUihlHyiEOrCSWh0pWs0YcebXy+s2Gvvcek78
fhkVxN7MyJawfXWdojghy9ifZEKbo0g1X7Z/lWlieZGrPFsstM/h3vMoZFggNi+lEm81zli8O5ro
KABEoeaVNohipxbGsZjazJSUOXKkJFVnElQUnVbj6oNYgQQCBbPnwD1SzqRZDW/GKW0t+vGWHOtU
OmdxSu9Bi+Ly//ssJlQIqYYmQ1QZdtALeLobSxs6iBdMtnKPVSs8dKtUx/PqKeOXp/RpCRVpKaJg
XHidKsFyNbr0p3LVu7gk9usRDG+D5MlLrlJhT7mSPYRqobNJll3IL6deGsG+cDaucqfN1IovFSQd
kxhTk3hIUc9N7tJ5SLWOFGdJNEHUbZx2zBc3WH85o3Fe/SJHN+CA8sweTUXBNhMHp6NsY24v7HQz
Utxloh6hsSiyqwNxq9s/l0NYBqqSJ5oHG3Vm1FhqCZB0mB32y9W1s6q/dO863UuaDRTyKsnR/vU5
N8kAasPb6lUzdf8qZsoBesJuThAcUqS09gDOtpqZfDOBqFlcZdZ/Mdl1gJubvEozHy0eo7ezhAPN
N3uR2Yr2wI2kxr7kd68UTeeAuQJWA+FdIG7GkaO05qh6pj8s8U35ongB+IeVczTkmkc++pj+2g2Q
OJAT7h2LCOSsjvLwqwpMmLedb9TX2teMJKMj63tRht1oFvX7FqOfNOP+JAz4/4J6bx1Sw+Wv+ChP
mh/s5GU9X99s1NC3rzaW3muWGrcUZBeh2LflWa877ReMx9aRnqjINWOd87cuto0PwkVJ/GokCtH1
nK55Yuwz5AIUxEUAh3JBka3bj7TENFDi6WuPbWVpZinq5cyMVgG2jE4UfzT+H0IJbK7/9y4RCzHq
3uHD5PLJq6OJcozyXwSUoJ8Ibg4GdRTD+/DTQNAt+8FVu5rpzs2zu6gZGMSGVdsAAdaVrkGv8DxH
NGtB4mOx9T3xzCNXGoTtZ6h4ewIN+0dkQ3x8UlyQG6TeyBtLs1Fon8KOaWoesMUlAtqd6DYQ6Ljo
k/KgwVMFxzjfWpYwZBeiR+X9EVTQOa+sqQDXOX0So0RXoOp3KLvGCI6ZDIYAkSPDH1u7J7mTMXFx
a3eo0RXc+mUviaNlJDb59U77TpfSt6x4srnTS3lzIImF8BAi9Cbrd/JoSdwnjDQSdiyxMnEiU2W8
f5vzIOaczm4k4hYJv426dpAi2/LOlJuqHqpyjUNGWOrKWnPde8QWpkJ875fzdmI14kRPowhxyDuM
Z8vF4sfPEh/DzHSd92iHBYueihYkFFfohDAfideYacM3ZevJhlmLSRU8MYxH2WvM8/kdWeocNoQm
ERPoykKP0wtTcucBNzse8yyWEHSXIX5XpAkU58yNdsU08slW1J9/VxkTQE+FZOGSpB0/y5FEZfr4
lwLRq+KG7MY328MP7n95Anqlf9FK7/ykF6cMGFWvAiXTTB9uwbdmubm5mfysoDPZgE056phH8y7g
Lvlm3P0Cq3IcKr5E/YJ2GWujpo9lnV4nHTFMV9hfLJK5M0qLFRotnLuEvbY7x2BKXOp9CUStIe5b
qNPn2WqbEgJzdyXvHWyfz1CAycIG5vRWcIFKmwHwRPmihD2JUHCXK3cQbfdtTpbAb+Yrg/V5k1/B
U89BK2fE1ymCG9FsEGlIgtd1AMScA+KHEo5Pp/WmZUVmHx85eUUdDDZyw5MxdlhEhRCGKZwh4T4l
jxZpEAUtRFRhJ2UdoDLnMdgJeiPW6O5uVkn2QzPLq1/m6TCjzjaxF2Ya/aoEjVjzDEij7kHnsUwx
xXeorxJ3wPlyu1gFT9sWdfYqTJ0ZbHdIYVJHitECib/KU0tT6XF8IDcmBpI9HtwdBjT2yUdeHo8J
H06j0Wthn67Hl4HRCuSAWmrZuAi8AM/3wBPZmFzMAWUUyLR/4Z2jqu44e9BcxthUa0dAYXP3u5EA
bn0kgbBMEAYqWBYwU1Q9w2Nn0QSr2epNhHRBFSoWFYDu3W92zmgPiGXhN3SfGsMXbwLHmUZaoe0L
M7h9tSd710+wcvQNQg4jsmrR164hP3mp0jf6bAKLIxkj0WM1QW6IOV/UXghrV/vrpXYe8pN95CUJ
nCIxJPLXcyv7gUYezgziyqSCh5aqIMJ4TtwVB+DR0K80dhjo2ZvjjI0M57EdBeuYcbcNBJromECl
tDw0I40qxpiUHkAzvFjCHQqMVUjttlU8yB74i6/pwSCE1/t93lzsXVN2RUL20jrWaIJ8dodwCRnV
oMMI01KZQLsGuOOtBNOyzYPC6oP7yTTHIHrDveG5enhh25OL8YcwTtW/LlHrn0koq92lZKmMerhV
T07vR4FrpL8Iu5Vay4KAk+8HPIRKkw7fuYncLVrW/fk7iNqR5yAOWqhPoTHXaFez0uIn2VdNNSFa
bycv2du2iragsnBLHIVI6UD0UMRxIlrMPZuVHab1utnZZ9Zce3lagIxnmy86kP0kadTE5AbNsKXr
CNlt1sYQbyHnqbrnaGEoDXBNisQvyLtK4aOxSxqJfLmjDz9WDkiD4SsqR2d5cETyPyWTifQtWBvD
Mr2LNN/1eawrdnMt0ZonDHl0wIqKrvspN9FCPqHIqMh981HTFd5NWx7He/vUGKgKeLUGY3fY0lWJ
ATN4+hfwgtxKptZvYNLYe8Tq10UL5sQw1gc36m2Ho+vVjgVI5A+jYP+zM2TRE3zPCNw+c/xd48fN
EwlXGCxwSdh6Jb59SnZHLIt9AZlwiw6Vf0V1BD4XhTe7B3XGcJhOq/MvpTlp4Peys4EUwukUYrqi
1LSDEmm3Z2XB7qQCImya219vgCNClY+qeV3iCd6iFvhX4eV58jhMobzY85q2A/y3I0LZqT6i+1e4
IuQe0Dl67HC+015HbWWWMPSeh4s9sGIG3WtMPbUhoIWXjw404JelO6suoG1QFRd/VKW17Q4woDZW
Ucg7fiLLZKknY+k4VqYAqURenzlee5WbiXcdSQ8vW5Pibjyc0jVkijox3zokyb7d7iWQFOmQH5wX
J/pRWRE4T/h0V6QVRTQ418KjS4EqhfbR4j1ObfKwuncN/nNGT5ayEdnDXLwBFtZv465oESFhB9HW
N9is+tv+m/utBqZZ7TOKp17HCXBQ/PlZqm2bHyyZxmpxIGxKZ16TwAD0gVbO+ZhbG2hJYuteXhsK
Sn1f8jVTN+VatO3ARdhkLsRhXeN8Io1B+YnKMTSfodvsr1s8IJZxpE613fvB/kUEQVW1+Ch8ZhTI
cjHu05Hgl81Zi/D7gchx9k/VFsujofhiiKumX2qdEz2p+dSi+0MiOd2db+C+qRDFBXTZzTm14JnS
aqkOdzWNfqjPU5xPlXNr+7mwifqOncRUYcVrSX6KaG90yFElHxbYFyJfpYkW+iPq4QC0bL8bZMap
Aqt6KK9V2GUsKCCsJaZmxWpKwQHO1gCPrYCcMMGA8W7JV0WWjV9D24SEucPEwo9MXsXijwQbjdsM
cG7QcWnohpY6R2iPHVkdOs8CI6eqa1lS73X4ZPnA6bKPVX4AO4pSxvazAA8UNNVGxa9DN/cQHM/e
yo6iIqXkiMhqPe1tOhp3etv/2ufHLD5EM9TByducuBHJQC2FssS9lKJup+7DVUPeT+fmHxKgVItk
fUcwjtKaSFP0qV7y4iKIYRCZxTSxA1x4psgRfsVF+XBRt7DDjwBH40EMiPa86FPWydCSyvvuixnk
pw75laGlrB39ZoqUvkBDFYDMkx03QgHIH9hcCsRuWSnxDc24pojqiidDthXNvTkFR/5D3XIpapL9
knEHl7Awyatq2kCjvVpFcqoBesO5yJ3rhA2XOjl2Ka4eNaOijHN3ZGBHycX9WifDk0lpbPrsnJim
PhqIyY6BI67O+15LA3Cntu20WKH1NDaebnq9obBtOzYHFavPDR4S0mlxnBPUT67uHslcFzBYPT3A
sJcKwcYd/QV3mlYKJ3PO0+EWqo2Zeoiq1nmf4YDVgpvPgD4fy/byoIRd4uJK0nvLYZvcS2DPSvOe
uusnq1mPLI6ez+kugXy372og8CeyEWjHHEG0NB03K+1y89xIWdduFcY5zJYc+5k1FthRSJQ9tzQY
xqihA7TWRXdcb8WkhGb/N3VMEblLM593HjL1Wqeq+UIhYTl+wErWCg9Cc22Zz73xz75fkSMpXYfl
tukXweuKmckkXMunHBT6eVPx2mdCF0c2iopcE2Yip+jVxNFli7tDcbmDSWH4rF3HUIT0FWUXr0by
a0XNoaXZCUi0tpJynTcoNc4Hp0Iur5mFWEQb2hjirR5g10uy+g9arG+UY135T3SrRQyXV3YgydqW
rp8cip518KQP0BYUsREVCxJUVoNsLAHHJHTELB1fn4dh95S/IiQSj9nn60imPCfsHszC8kcFwqW2
hABhRp3Nd4rZV8FxjjzK2kPx1ZJySuBmkTC4IxQEo/8f76Z1+TNbVNf4wxMZxuepqcAaQYzxAD7n
jIDw7RWY4KpY3dVDxX+2V4MZFePooR6dW5pFPu6uFQ7bxpYaRIE9qtzmDRLUS0Q4lLy4ulYe2bPT
19zhm4Bj5vXX5wt4qVEiCUVlvwGWIOYTABwoTaaEhrji5OgliVa9IAtI5e5YwFHFKjZjE434lSU4
oPNLsrPAsReTj043zdhrglqjh1aIEw+w5hQ/LDXQb00X6lkn47NZnkuVBOvppnBrWeAjwe4Kawpx
tbz2UgAhFkknFBCjXjrht8ps9z3EhJCp26t9rcq2tUOg2AVCmXdqb2W9wzUTrTCsZUKUsCfFObwd
t78uJW3HKxkaBas7O9KU5BeSVRDdLgK42fzrSEkp+pYIO9KJ1rjCjjDz+xOjgxA5goSiaxRfwgS9
p9QrYGUWAZNhRn02DTbNqsk+LhrtHHJMw/t3NBS77rvudPp4/YDQAJOMWvupus8yNWPhEo6W6WK1
ad8U5Gw35LK5aZxAvIq5FjxNxmCDfiVQw1M33jUi1UtIMfM+ykykq9w5x3i9v4qWgwUInmyxGAUu
3bfxzEM/9Z1houPVpJXufiROA0A8vkFzCq0qaDt/bvwu+AG5dfhqnFjKAHXY+El92raYvtmyjfm4
HY6K8nfEmRB0VS0BVJScQV0spnp+x5P+7aOJFu6pu3Uxp733OkPlNE8n9y6OttD2UCb7SMwO7zlR
haMlJAKrY2lU5iH5zhNymKQOEwrYfT4SzAa9s7eaHQPm3WOIjuTbl18ZUnghLXWsKPA8PSZrKCQQ
JMbLUVBCBcTguLoIifgACouEA8dGs+3jMo8AShdGx7uod/UUv3btDaBSb0uPJH6fIGMthpypOvnL
s0ASbvjpJsbSz5ifZX3cWZ+G63ieCTd7ki05awMW5qtYwKMX6VfUoKjhAa//bix90j2KZTZXQSs9
Pf6FQ0M2xT0hyqYcFMjQodzIrMuKxqBg8bYmhRezXDxx498UHuIXhy32Dn2qaEx42pHtQ1cAiwX8
F8cPUw7PeebWtGVW0TALrs9LxxP7iico9RS9p2x48whKGOqnfCHVWv3HSG3lynbqPgQrhce7XaEb
zc/rE6+ouZDMIL5piKc5+AqHuYgYOgwYOXg+fCMyn7dRiPOtXQufQoUEHeY4n40Haxua9B4B9d4N
k+nn+rQRuGKdBBiASn8fqLyCHAhZ2E41/BfSQPlbqa6UXWaEvr7Ob+eoDhY1tIjHrq4E0O+tWyqU
xTQuSAK6I2TSDjEcJIsUmzsa4bcQXtfBUiPhfzbV4FJDx8pJxLickPSnVZFmHOAbWmNA0qgmVWX2
YkN+vFMn15v0PUUW/6T1ZaI2qNjVlN35D/2Dy5Req95ESwRudVE0K4bmG2IZK+GvbrmZS2jfyC5z
pWSCbNtMmkfXsMTr0m80Qh88mvAfXzyz3qEuS+wnsR451LiuS1r8KUpJ2pYXAU5nx7klKobKXL+x
sooGhO1zHJrsvrtwQhmEZBaodRK3NsgLb4MfDHnTexPs34+2qR6AVc8iqUjO6672FDCjTjaxdH8H
H9sWMhBK0oH40JGsrzq11XzaU3ZnQHGLe6iHK/yAmtDdHHOAQT/oj6afHPgcT8cO1y42PV3zBmUk
vFn7bWe6087+M/KQN/ydZWGyhx2ns7O2AhTH6wxVFofGOmeaPfSzASvAKog5HEnsOiyze/Vu74pt
tV/HEfTsTfJ1HsjjL0trhJ4SRCb1j1w3hfI6TQpnZjmKFZJCc5QB8v75ayQ4TMzKwya9roUHxcKf
hiklco0KVFqgMcyWiTwrJqNSvaOI/8FFhVpJUM2RUc7Yl9X1ktmZuFoeO9xWqKOFlOMUWYLm25aB
vO9BZMjQflXjqSf5/OsvK2dIvfqAKcWBSjd9PlSbRllvIzWM/vvsa3eMMBrWQA+vKjULOkT3cdbf
aNYmnM6YDKdkN/EOJH6WjRKv5ELTFjE526ajdfewrS/BZLfe05reftm5QzInhWfRfsENGkdvJ9oE
ieatA3PLj+GbHoUiDqxap0ztYcHnMh6Pk1suZGsFUAtqKYC7AEhSz1kPnLwIUWT+Kogu57qJ9ZJn
N6Wbhqq1V3VzXkYCkAL+3fkC9IT/3z6MxA+OlYwgsyMfsQVdt5lXDbT/krICuv5Hbv4/v5ACUplV
GXPWXMvR8zuhZfqTaghTHyodAMfGdWqQ8I0XafGdSq5Y+XbnzGS4bv6wE3J5aAX3G9yq7+QnVJ2Q
OnBMhG5PhHmTlCzExJEBKjbI/KSlyWEOWLlLZ2CIViHqHQ9eIG2QoPtZgQPYbBbdtWQ+Taor6CPJ
onUTzAFPuOaighb8oMBelXFjyRDLz2iu33Po0OUlwXPIIN3CGQsSWRplyZR4tZ3kRPNUs2z7VZPF
I94oQyJ9NzwNCVlySCfm94MSpe12VXoSeHjmKgcsQ3bi/KghME6nIA17/8D+f3sB+V0DuMOUoCEo
de6QqDelofVgVHi/TrwFdgiP0GRGhA2hhS17g5Pbfdo4oDSdUU2ZxoaD7nH2mvX5ZR6JzG7uX2k6
gg1e3zlQqM2xKWtEKjz34tYFQHVeofVH4gVU+b0Y3+cgaLpjil+ktfSs6tuQEte94aPBvi59OCtB
QmJnm0CI07o8WDSE0Lm/3/e+VDLg6ieEBz0fbGXyvo6PonYu5AsPvAmJC0vmn69Vq0QbE3Qwk/nI
7+kcmviOmHZgqk2bxCS+hiiN8hwhUKTvirqh0pj/Y8JR5cqgoRSE4Rk7VlKonhfNwVOs/ZR+N8C2
rHimgeS5qkg4w34NDFvLtu6Tz9yHsbHR6BPpqbJsaMK40LtgS8cMKVP4bzUL9tCm++0bOwJEAXrj
I9zloOTIFrm7wcdJLprVQ94EDBJVJp8WXQIBnvlPQrhIwcAbMzqHpHZrHn/Jv7dOwarcUPaZ+vXy
mzSKi+TzElffrPCuRTLeWni+NdFvLK8dpdv3ex6ncJX11H+pufxX+CkbmS65DcZ866s79C94Tr/0
QXUTNfKWoJ9d+QW2PCIEWi5e0E+l22C1leV3Xuue4DrwJnedaAjk185WCNxNsBP6n5cR8A6yzasl
qLHQj+pukCZWoG8QUuq5Fl7R5pSgiTLMYO11ovlub5pqkrV5loAfrIrwBUeT3NYza398At2qO9HK
mSn+YLu6JQCq5h4kTr9mfY7IuoiabG9o+DX249xT6sNhZQ3Lhrfw1jDNw8ihDlmGvQVm1WbC7/Dw
A6kp2zeZu0PqhrIpO7tiEwmufxdOgCbr8Z0x0y81jX273O6NiWEzlIa2ld8H63Pwzx5MJ1LUaPUk
O+4xhsx+7BClCyhP6xPjfJfHFUBxXWeqS69KdcCvNQ8BnIq6x1XJAexjD+9iuGMtrG2ivBd3f6j5
zv5Aq97fV63cO7LtRQcoDyo0nuMZQjEyFPZXBLaifSRZXULoyKiZz0GGVx5cD1GNlAp4OnTjd0b2
JpnlPkkzK3PWaN0KDtJC4EAwNC34TJFw0LeAcFis2P/qiNhicckoOCloL6Wkp34eMRqLxKN/eAex
X66IW9ceMYh5epCHL4SxShiumvUpgfhc8FKQbOMtX7Z/scQCWOOaYdB2LsJMT0HzgL++oNHrNXHl
321oS2r/aF0Osdgi50sN9RvKKlFu9EVyX93IY5sBdX7k7LwoYpaQ8A2IzjeUaUYuvZGaNjsyVEWr
1k0xZfduFBvj1fVwoVk9Ic5tpofsd+/XIXpUYVfeYkyExWxWCCL5P7EqqtvO4EfahTkdI7RJgKLN
3jsjU7xgzbUfp0Ewk4rLxum/b9EJdfLPSE+Sm0FQFJGRrXfvM39v4AqiteIIiTqse6SdK/ASFoHG
PoHY6+unsG59NlrHAAhdSyUQzc8jIjtV1v5VUDbOMnnZcj1T2xVQhr6Yti8s0O1OSfxDwrF+QMXw
CGu82DYt7VucoypI0DwjAb5bf7Ex9q0JzheHYlTHPQx5j+I3MIs8us/bl+FDhjFAvSyX07G60NYd
bM0dI4LvrWAQHG3oCrYSceeEdPi0b8UouTqstbIbGX76XhFNw2D4XElidVqRiRN5roq3nRZMMcSV
c6POeoUsCBVx5LA3FVJM0d1QM1GmopEPR0gFYxxACSlJW4MFV0G4Ga25fYmKCRiSHC6OFbi0yetA
5vQVWBWrkNz7sl4ECt9BQKnh6iNF7bBSI5jG6m85jkj1+9x7vx9PSPDY06TZXMaqemjQBCPKEEEg
JBdY+wEZ+vUftl33WsnmxmL6LAUFB+Xu4hmGwldmpIYw+DyR2KH0E9h5ZL5k4ruc27C3ZwcS8t6s
3UpZ6kd1Ose8/Z5ibVkM7WbzzvylD3WHMIYae9JOTlCLk6emSuf6mB3Z5losTpFx/KEO69iWNDAM
iDMeHVQDk/kUcCe9hllt4QvrhsqiDHTJawgOpc7139pivyLiSxxApn3o7/E7sH5AF4gDVqem2GT2
Ps0WF5joSSZbKSmZy7+fijPiWqS4Hg9Ix7j07OVoqapJkyIhmjmDR7BrnNhE/veY1ZfPdijfZecJ
CLc0Zdvd9oo7EZl266JKUYetUp60Z6qWP829m2fS93L9Z/QtDGRdnXQ7HhIqD4rx8zBZl5LqjNPC
svoGaf9zyMRQNNzctCmeProaiLyRwH69zDAUlSX6mOVqPqZoRggDdwDLKA84SfEyo6mTILo8xG5k
7eUrzDqJpdZcv+HgVl+56s4jQQd70k+iUFPojTBTHF3F262URxFQIX4Ja89tBgOYL9IT1NTsJ9IH
okNAvDBcZ0kI+dv2UjOyg3MaU8orP5eVvCXnoSD4fSIj9y78AYHPef8CNnVpn5Lx7KA5qUScRtel
58yXJD4j7Y3Mkn/+h8RsjUj5doxQ55wKHLog7XEV2pVntQdcaKLGN5neds0PnIAethpH9r+ln6ZL
gEEdIoEeUSJwfgv+VQx01ytLB6qax95UQwXRaFjMk6oHC0MSN6BNvSVSS4fQnFOO7pD0i81vgo/F
D9roBgYeIj8U3Caz2UkMY3Q9sJ7mbfV9iAm5yWQMh5pZ9jeXXatXWYlnv3sKHrUmflYBDxB/u7Jv
OoNWWVBpCzqFJ3FMB8z2Ucor3lndGrImj5d9ZvqlyigaAnxfSZCt8iG4pdrYZG++7cuwlUoS9upE
KAQd2q5GEvuKup+QhNENpsN4Eo1PbMz0cA7NNk92JJuCnT2D5y4kQujC1hS80kw43d9WiN5EFrq6
X7+snBSjLbThnH9RBKjbI966K6QKSg1CQ6tb8+Xaj0EfcK6uJRAQ7695ZKMYOYai/cInHQQao80i
wPh9l8GjG9ckcrpK8Bq6RrERktU4OCxAtA6Hpvx8qMPRWTaiN4e+P34WqGRb0EZYGmjOrrPisVpy
ofNNTFSPSmNN3hzRNNL3bQ9XltCkOdyNkkAH0rluJxJdRl271TaMbyz2SB2/dSs0HwEGYublNEG9
8oeLvfv18B4l6bm1ElQYp9mC/d++ChBid8FDkYd2UX7X08i5Ujj62Imp+omAOyhPEN4UGFKIi1oS
FMv1b5Ekkl7b5ab8UB7vWpnHFAhnSyx7TgXiyqHp6RAP7vnC5CUXms1MW+/Dyfct2WV2g+S3QRGm
tvvd2dtj/TSYrw1WVMM2S6m8JND0Zd7vqWVkpeDvMRIBl+XTGCMUZaCoHYM3TeillX3Dg+jg29V5
chkkyj9vmyTH7JCO0bPxgNDtq8ISY0TUeLx1yI11Px5AuwoMIa31ANfgCzVHoHTFTIgZdHhLXmtW
ZVQqQNYJsRu8QJOlfpjNLe7ZoEZFB1NXsa3PDENya962BfZYs1cRBUUjc/CFL0XakL4NbXpNFCWg
gXz22WEMgfP4Tm/j3YaqVC6ue3n2W/eJBj0vq739EmVbOqOfBnM9XiGgwEtaE0rmIdu4B66akJ63
mFyD05St4hNquK8QHuyAMkdukGidSTaoWKNpkaC6JKe0r1Xo28wNinE3jnAmhTJoTkKoFFpJsUtw
yoMtRO9nfI2aj2JicXSgZqNwSOmcprBWsFNSRIgMcpwZKLP98U+iZTLFe9fp5He8f/6OCqRnnAIL
Qu+8Y42uYAYAtMgnc60x0sDW+8GvFxJcfpCxiwial3OR1s02T4Ah1qD2TZoW9+dc44OlqitdE8Gg
3N6RB3j6JSh97IH1NmnQQMR3/0RWqroPTtN1ufF2Lz2vg1NZnB4nv3f+6Hd66d4kl6NKz1dBV4PY
Q46+spSCbNHFTO9iE+uw9WxXkOir1cE5kMwU0R0vnnmTOx5JFlu2OqnCJIzUOjJkuS2A7FW3SW7e
KLIFXfg62R/muLqtdUkcnZG8IKh1TBQFrUUQQlU1DCMq8O+uWaNGfpLQCXtvOuZeQ9fyPWlZ4hCJ
S93L//YY134M4QdjaJ5ZBq/a1u609w5I/CdSsAC0h735QV40JgyM9bH0tz1A+YLuLnVO7BOEsarR
2gTLHqfqsE32wPsURlPXS2lNwvYGMzz/lJFo2RPg3uXaih8/jRlhMHMPIihhcNg8rZZqoad1/NO0
cYLvABuurM8QUsuL21S0NX0aZYe2JYyedCrpK7cyxtcX91rM+hblOyaXTenGucfKljxf13+EtIPQ
IGWFAV4R7q5m+FK67sLPnZiCq9CDzz4TlB2dHfo08/Q7ofKKmFiEbS/YbsMF1P55A4S0lH9It6nm
WHY7f+3IYXN52yOIjeCC7ySMuik3xPXPIHoiNuUt8YvveJ3EBesTPSFx3ApO6Mj1a+WCS6o3aSIa
86kGIehS+kgvewpN8dHpf7dHDdvLLtV5bilJ7qhHUAi1xDwPq8Ec36NMXO6T+aSe9CQ5TMVHX5a5
hFjDQf5MOffaHFuv4eKRHo306SHpeM7qnOudYmvfRhFcP/gYfKYITpzU+E1N4l6BjshPlY77mXFk
rLkURJXMejeoOR2zJ7S/JPEp+yOCGEmxSmAgD3FkH0RHpf4gHnqwLsXDJGsyXmogboFQuXm8RIRR
3WiMXzB8J/fgyo6LQiQ8XNB8B3KJjAuMvgndXFF6Gxag1OCQgiZlOdTxU5CO462w8OZVvL2VXAx5
aDRW6qqyqra5J8ISfiLvTvc1k1Vya4dHgmUIoWPLwt+PcKEWhJ/lnwgxYuFX6kjfr+3moG2z++Tn
AsvmKly/LQHvIsbOFwI1gvKzT+gSmSbPnwvaZbxbVeCinHnywT+PrlC5f/p4AW0LTaY10EE9Qpzd
8aoCWQkd6FpEXwUQd3EMQHkepXxxFTyQfqDb68B9A1Ep6TSZpPYNtOpUiN3+dSWK21OMCyTckS8E
5VgRtmB2ZZsA3qzSmjWOoDtQRbfl4GtLwqYQuhsF8a05tuoWTFG3XA8Wh9K+M6Xhbyfmk+nnAj7y
xbq/hspSnZHZsNVFlIW9C9zH0ECFJLj3a2NATGZXObmUyV6XufCFwkLE84A0rW3g2+D4o3G7qoBQ
ZODVACCx5g0aVkWhyLLYzWhTzTbBLuWZmfaeoeCuPTmVQ/F5ArOIJDMbIpG2wyD4gk6X6BQ/ZOtt
FCLgmdI7Sb+vTIo//FFrUGMRxgfKDb4p3uRPZUNK1TryNWrk2TCYCOJbjI2bAjaLAWRzSSc9Bs0F
lFfVB3dtcyjPPxwbiWYNMmz0fSoNBtnZKzVi51q717BmIlaPUqg77tXf36lfIP4oJI1Fozz+DyUh
6AIi6cXJrkonGLK/AjFjBeWsUKpIJM0sMhPaxJfffOa8/5XrPhFi4E0jzuT2AXshrPnGVQc6w/f2
DCJpLMLpiUphzlRf/1UkPDJztBYpomZpmUizKG7wZVxcZCpkcpKlL/QkMWtl4rGKNp/DwUbk4vM4
ZyzbDzhL6acQkiUIB4Njke59IXtlp0NzVt+eCupNlHbcqSxSYsgMa8eYnObqOqiOyuveZh4+LlMQ
tMReOQ/u8rqWRI285AqfH6ehHFVi6E6ZfUqUQ0l//2auSBlb5cEEpqjFRZjM6EJcyTsErEcdR9MM
xuST9BtcwdOZ2mZ2/X8lH73os1lClxZU6+MRUXmB81bYpSjQs+kNueqOm1Enua0UTlz25Q3M9IH4
08d2QVPxdiFC0pAygHZ4zdacoDSFPMGEyeCydk4BoQmZt9O4v+cKwoAwsHW8BCgiOlUrKJfUxQSD
yRdGIBn+kSPm6AX9RFJSiIlpgGVC1yDxbbmFe+/M1h5Ckc7Ezn5w8urlfA5vcOofCQpwwuyMyueV
r6YtlyJpAyKAdVwlv3veLxc3y4oNI9gi23/usgxlVY/eHKIWPVeDfbM7Ctoo9VrHPUlbpZxXxQI6
1PZ3I3Blj6xyHTmZzNl9hRYwW3mx3zt9eQSZZBQijc4te+yLdD1sZq2UPqqT6CyZ++O5JxPA+8HT
n74rO5YC2nk0dtiottqm5uAvRTC+XIMQSgksBhy/p/TbkZiMXgcs8tTtH4fQJ6I2xrCvMSY6R3Fo
6GD48uiDjT61uOpWhB3USR6dz8qKWI/Cy+vePKCXfXzBfBqHnhT4BKfVC0S/AOiB8Mws7ctbo3PJ
XUpB3vgUBVZP9fAmMzEkIAmgGWeZ+jBFAoNFo5teRPkhDBfmTxX+yivirbJjhdwbVcNRTLtlxJHy
zZVvyTRr4iOxJtpGmjKWc6LLwZk35vakslNwTK02w2XmNNx39rI7g7f7KQ1Bhl2IkmN4e3uXBv0k
Rky5G8HY7/mJdCcTnek6oz47rsj+SekIlt0Y164KGDkxnZG79p8/ul13QNSPJwLBgeNZCs473dzX
uDfEtBt27vmDqeU8rDfKDuwKiZyvnUw+RyeXY/11+w9EKJvBAf0HtBAxfBA35LzxAhdh54nw+/gR
he+sGQKLRIMqd0EpDC+wzGbDqxylOImcMH/kTNmWOs8LKVdjNmHhDuJSjshyyGJKxxm132rocXSN
ZeLyxxpD5m109E4gCkhyYqYGi/iyUTn8TXtCgTPm7oeK5D0ZfzLnQVYZFUtBf6usSWFvkN7f4VrQ
Z6I0sG0Un4hU3Jfp0OWT0BTrnja71Vw0p7GleBPslcko7HLoZy63eMd/jFUV0n5lJK2WYmIoVmdh
uGlQKp7GVaCE8emyTcIQ5zaYh69iGaWWo37slg5y7rePsEjLOuzS8QKVvlFiydhcqKVnqpMDP9eO
sR/ut1t7go5c/lm9rqH2ulVS/+aMeG3r6Dunozydu+DXcjThCeklmHi4g+pj1g/2MfRh+tMbM4oH
bNxVhOf7gjm70aLsWIrwel71DjF7omZeGQKB4YUlKS5gESJ3sEOgcNI79SHC8vc21DUZCuMfi/JJ
ZY032NP78C/FBmzgLPihP+qP8DJZ0ri6utBGMQ5Oy3YLJYoHK2CpiEcy5fj/0wIaH/p9UWMw+PJG
YTQ1xom5bSlnIsRb1KdI4AAHI+0tIuBRDAH8yapErUuYxRAe6yZZIX9oLAChrSjgg76QwwfjnwF4
WCE2+OzMd8rrI6qycrvh2xWaPZbBUKfWGQ9Ujl0VYH84E5J8OXiLxL4JwsjDazu2ukfRHus8zrtD
fxYnpAVIe2jg85/lzLExBRaPQ6IQz/XNC5OgK0zadols1qTVNmpq2nYIJ90wm1bQRfHYP59Odgme
zfktPUeqGKxmGhYS+BwghCItxiksXL9CaDATIl2mV2TYvNJpHpv7Ma8Ko830kiLUxK6BaFvf5JN5
L77MPWmUZ6FBGDlO9HC81HU1mY6vd+q37Ai0XWZSNfv2qymNJndm1DJQsp4Mose0dfah0wMrdacP
h8cT77SWT1tt050vo5M1r02QlM7/fA2f+9OqsgIwaQa6zRAn68frHbaFf7paEFnxkvqPkixh/WNb
07JpCBPWPQCdjTY1UXPa3NS4x6s6BfQfed3jySrmeagFMZ2QpSgGiLNj9n1rB748sOG7et4OqJSb
2XbIGNESbvgEmiidYzrdkRkdpv5yQGVXirkJJfRHqjfj7owhuBiCSASgwyKv3+xHDgB8fgDBKYbe
tzCDylWgsuLqhDuBqSSAApj/CrmUJmySM2cQdKLqlxGbAWjzjApsXok/YPL8MoqR+7gT86VfJZG8
5A9UW+MIPW4DhVtYrLEbT6r7kFGh5jCZwEQhsKt0oaSb9gn+dx7EdJjxJEQVmtXMretaj/n1cODg
3PCT2sb/ES5Gd2tjRe2Z/52tET1pQ8q61HgTsetrCyqEr3yQjmijSBXgCMoRGpfGRqqTIjtRsCFr
r2JtbXo9o/vXWSkT2pST/4LJek17t7m4Jx0F9oPTn1ariikoHsndfIvKa5l5CNM4rrAGFP3lSM8c
oSmGGhK692Lxt8arkTZCBrlyYn6RrDJch1N1WuWqnJ4X6gIj0QgDaS+qrNdBBJ2pwrCcbptZQ0CZ
sYtV+6dlgBEc7ZHIWDcLunZOuhxT+hYf9TO3pSHNcDVSbTs1uHU4kk7RDheM/4IMbjdJHCOnlcQT
2IlvzSOkVQTTIbKF/fQgQO8C87jw8l7Dtg2erEyuuCN1+ckAMa6bkuDmn8vqfCkcPpC2CRmtK+4U
vKulyTDV1FGg6BdsLs0NeiLeTsVRju9Q4Z1gCuwKE80Ruj1++mzXJZiP7h5ANTyzjM567OcRXqHV
pi2Iov1BVTK7U5pRTeKwjl0JknxlbiFj0ihtFbnyTToBOyXbWI/+2j/nj+9fuK2JnYdr/CUKdVBC
2SegVIbYda76GQoal2R4NWbXWXMEwSN8xOUGtv2ykAB3Js9uiNhwJI9o14neSen8c8GY5DX7dJ8S
NM8lgqYZvlad3mbaiVfcytCyo4C8Bgy23GzyRJcA5b+e8R6cfn4U660jVfRTCOgZoXDQC0XIzao9
dEOTaXZj/ZGd06Yd9Dt8vh4pAVhiZtAXdv6+iVWe11nnQq9FBlTV0NT9D4cbAkY50YuYn+FgbIoX
6JmCmNRAbf9QhC42nNMJSjtn3ekrj7uA+mZEdIEL635PjO5udtYfIIxxw237UJHIiTU7z/FFB7si
PcJth4/It6x52h2/sS7Gze4n7bB9rDH5cvumn1AcuFAdOP6afAkSeHlg6QMSFuNZ+q2eIJ7sfl5w
uEuDvh39aktUeBEfpzER3wrASiFsKhjI6vhitNLurbfrM1a9S7BPioqaQCdBWV/Nab2vWWWZ4ovz
kVt5IF8u/MSMBuQYvfxmL/tS3BUCD/C4wPf5a2CZ++CPGOZ7APfzhDRUu9FtfWWBzePGuScWsMjq
WbOg/y5HMQAKiLlAXc3jQeYm9MI0xCqfDOuiZuCy/f0V0BspOtikxBHcRumHXem340ko3mYIOOdO
Min7LM5BcNZlMy2nGX0aTTXiQjgoQuZbnsLHeOqoRoc/2bn9OPvLQGBLezpraqymw29Ph2A1BnSe
SFpl7EA4GrD+IEdF/DEQ2I0vbaTdeB/wfpT2RRXTsPbt8AuZH4fDxcXHUMvRuxm5VsMuonYJ4plb
1uCz+lRci6kxHxlMbvE2+K1NAkXZDpA2dqkvEf6TYvvcI2VcYMTK6v2aBPe1N2TOS2dPHfzqikLq
dqt7sjrbT2HSwG+TgaJ883SBiCtJJY7t4tnmMM2wV2/nCLLZKgpKzl8XlBwIk1GsRxHj2UZb7TPR
9VfyPupTLSv/O6KacBnZ28fiZAm2gH7l1GBZfX9t72cR5npCgowJxUEbDDCv6luOAq+19kcmysyR
uBBTswpxQ8ZiTjIaBI+EQN6J5uGWEqoBBfH72pi5u/0iB/wJ9jSID+dDvaPghQkA2F0j0kw016tU
Yntk51JqscBdLPmXCGWRZa7yl/rSYJXF8wl/Ti8rn2IFzzAgIiy82I3nEB91wmh4PGe8XUhFdTOx
IqKwCQN+Tf7iPZmEbq9N2YWa4VNKJgrNe4Zdw2Sa1Yho4ItxUTHkTClAsO5wdE7TjHaB8Kj92vR9
ieVwuZacAG16tZO/B5tHK2h9te24RkZ7EGIfVndMJtqvD432LdbW5pe886rEcE5/B3jm98Upd4X0
OJewReAWWbgThFH3vSqD+e/rE7l89XL+7XHXYd5uQopxx6DEymmIP2hK0h/1xbRvAlmQ6p6DpxMP
nnyjWpSbkJ68tvba0Kjg158hx89qcBt9oXryr8CX/w/lLawjlak6IAYLAxL5gQoyoQbLvO/zUPnJ
RedxzbcXFlUo27PN573O6HcJak4WGSv9QoFqJFMNur8RvXhPhYnBrediriD6PmYzcslBxpOk6H6h
XAuF3Yfx1g9oMNeosXljdJbfnwVOR5IaZ2mfhbMjostBZBjauJH/ajwj8PFTjfV9oTx4FrWsBXuj
UdE9sJQxUdLwXPyOpgkXPOtN91s2cbvAgwbcfOkg50EG9PUmQkBuHEj+8roKKusD7kRzGYVMrh3c
NfU833/y5UDaxRqgkvE7FBbkD7iRIVNzSl189Zzg/DN1FXwLQWVqqSq9+qgi74GhXUVBT9P4C1Uj
uH12agYLbt/G6LAMCWI30DPgIvAX7ZQN93aFyjDKBMnqKZHKVxPHL/qfQ5Emv2SvmWkXwS8SRI7J
4fhTbX6nGEORToQMxQ/LN1OIG34DHjtSRr+qcR8i2GduTcT90a7FeLyMKOYYuFihpnaDnKwmZgkz
i06SSFcAs1El+PuPIe+/MtLqG1RNGchRfVto0gEMRWZJPFr+yB/0aRLZQwnETqUdnDvXzGN6wCZC
eOh5fZ0DLzrmTAF3OB5asGnkhli8T/O9YYpPzyjA+iFIckS0g7fsEzm1mx9ZIq+aTszf0IyW8QcF
2Qo/L4EhxJam3aTWy0XMQ4yHIFu48fMf+jbKowVmvYG2GCPVvsX89VXgi4FY+vzCVl41LbQ594Sz
TGEsx5LaT6uwNKR+4qstMzANI8npCMtX4hlq24DYXx0UPaa3dIIHy1WAIGDnehKTVWEZ3rMzlxLv
qQBdcIRAuaLBOsVPwfakAQdTCdxMto1Sh/EV5tucOHU4EnSKm6bDialG31yHh5iIGEdjb7X6YnZo
QXHvFHhhJQvO0NAG+A+nU0dBxlUJ7F7gcbXZ3RktlS7nrBI1sZvHl8TmoKTdJmD9e0SxzAaXUiSM
n+V85WoeiM4FVEc4K/48ie9SwlPyHj0goHiCEIRrpx9tqSzqW5Rd2kWZzNhhZY/l7e3VjvihL2cQ
7MSz1sol1MUfLgInkf96XGeoHBZ3tm3zBKlU2FhPUZEJsOVU9ETaXqDy8GToRqbyKvbwHUOZ6QxA
LkrufY5RXRKmoW6sxaNmGcM2sc86ITsCk5c2vtHgDVLKr6gztA8geJbrzQJZf3360AlLt4aIv36Y
mBfmuHWpeixsdlEiFY0qMhLV10UEa8MpPuevGbLZIZOjdctaRlvG0WxgLR9A2LsQDRwz430bm4eQ
3bVqx/x8vl8mYdhXkdZyYZPbqw+42H7UHHF+OczeAK7jfKYl+0cHX66MF/SSu9oS8kSbgTiYS5ev
ClPYNiMqV9TnHCyXqIJEh8TOyYFaxEe10jFQ3MvODtVjM8TLM1V3SuL9cJgYkxZ2mv6Dms8aiGsO
o99t12sW5ISeQWZQy2rSxrUpOHArOtZ+L0Gi6JYDp/1Oy6tg4xh9Uzr7T0aHslvOSVlrye6fH6f+
MYjZ6gtNFtnFe2rrWciSHekWNOCxCYRXIPmMtpX0TOLnkBu8ieuXxiLU3R0ygJrA8qpwzMEn3I8l
3XQ6I0I7C1MfBG8jvClb/rPYDe8LnZu7jrdFy+vZVD5cWmKBttlP/g+lJlpTinHsF1SAkoCC5+f+
jjXB4LgYvL+VVwntHS71d1kr2SevMW+5h90s7VDihKy2Q6ZpdnV4Nj1dYoUih/SLKFMsueuXDsgB
IMGraU6j0HvIrGUK8S96n/4u/7QGxwlbLko7WFkiRC8GLXkY/RvxeNQZOc+LfuH91fYKgdDxj5vW
/Tal3XNuVYy/wf2uQ8SM426uuACXKBOzWW/y8dkFxGkLoKJ1A8eb1/thOdk9HqDgP8KE0fkBph7B
xKbuMdn4bKXmWEiACPBpmWK7zuLBtKYPgf1UqyMP+QY5+zgJNJ1YYTLwiP7VLSysQ+NVXJmoE5lg
YuD114xNKusS2f/lM5458OGidzF4iD3XCI5NqpvbBjK2Z6Z6mO3BV2fLL5HJSJSTygeSkuzqxImJ
hnDcHfHdTinu7CeMvld98x9t67Sel5TCOX3nRnIGMn706TGkPK+UBgHNwdMyP0I2EtLazvksSig5
zAI62aK4d8/K/V3OKEc7wpRPpickR0pgWqlNOsEwAH1kSwEbuznBdvvmRuiMZPumWgeQ7P9WDbUZ
85Euu9MC81e1tcqyJi98RHro2Uk7A4nF5hQhdH9MpFTjwhCAgR3fHJyKR9kcHvB88co1DN+DKVcr
+U2H06MkZtdXPH4cOnqCET2+eRGdIdlIjS4AW6zNGGH4hZqLNtO1rKevvwPthM6/3dNjSoom6D8s
ZD0fyC9FVk/iwnOrS06oJJejYZUwWYwN5TEYYa4/K0CHzXPksH1IB5JqMhY/S0a/Gn5Ps4V3ORtQ
X+ekSiVEhyNAmzITQx20ihbnDI2gxbX8L8h5iCu9Xi4oU+zmKOUqUn9m3vj7oo7yYqmfOr9w1LO5
87pvNiVLop6RfvjCr6Y/qA7vWEA3POjzZaccILDgLXcLYa8M/DeRyV9dNgG87bzR17g1EK22v+UY
60LIJdrl+/25F5hHie2wcS4RYkHSFdWSLMMn+gh9Cn3tP6QIGTCxl6EbmfS/jLGKGGIlQ8NOo/xE
deDzg16yEAvTar1rHjx+C5EywLKZs/xwWcagTwV92nUcDNIoDo7jPz0GAmk3EPUI+lXTOGs52PnK
2dXQMm2s/ioSdWdZODGHRGVOaXD9vwaY7igIatoaE+kq9gOsp9E4nmF8WMe2/lXQIPeA82t/AK44
pbo23YesmqJ/H19dk/vbYiL5EaQse7JUfC2uWriIFTFwl5uoJ1XdNMSpvZgOOpihggh87eEiXx3V
qc0vJABMKgt1JNPh+LA+oA2kVDLJ67QXJMpjs3HwRdivkm+eHWxpR1ccKcDsJwHdJSi2NACR4X2T
uGjBErGgA5nCBPH+ysRmJkczKx1XOU+oS6k8RBLJ30LuEBK0v/wvyjBmuijNNdPaimFzCVsjHlwa
wImK4upAH4dKg+cG+KDipi9EArjQtYrBa5CKnXoeSIQTG56tgR0Jp8p9BM6yeYM5egFvIEsu6Lag
FDc5ncjF1elcTJJakdgF5x3qdUFlRvKonnVsgE4l7uaxZSVhQImyMvfROzJzNrzIq8cYuCVSU3gK
oVSl63rkbwX8KtNw0zyqvU5ruB7NXBx0tF3iZeeUnjVdOsUFVs/NpSTJYWYl+6NVKEJNGJsOQ2n7
KXTw6qZt/szORfzjAzUCeiXDl6N1ePlLdsyVzkMDqhSVUu/8FVFHIRAnEXu26h5VNTg98vbCWMrj
B7XvDVIEUrCohVgXb7WeCHu9y23POGXjkMycXoqEtfQX7l2Etyb6e2jlBECRjXICXktOKQKX84Ra
2rEF17e/blwQle8/K1FkXgGUJZp7h5qoob2B+Q8mdstPARduXIpeamC2dcsGiw0gi14uCFcHmDo4
WBq6PVHanB+knu4ONkXx+hyMDvxn1nyH7izW8YNwLI1KYhr7yTVgkGr5/MYOJNT6zCeOkurKhCy1
VaPuENWeYLdYL7NZ9aFghe66hhAy3kbkzjsB64pGWZYrBWJ6CszpajK17MZn2E+owjWeHx9wOudb
Ea9py7gXcr8aMVJKLnLidaCbMqt8BZtrVQsc5iyxCmn+JJvWo6pBJjwlbUgakENg8YfLMXr5khaY
dkyG+/d8WQoFhc1rRQZ2wGcKOLgmmIukZLORUumVGUO5oZ3Og2p3E+uopgbQRz48Fu/k3TpA7OgC
dCCgUO5ICqnPs7yfZTD3SXOP8UiH07+6qj4GDBX5S/ID+nrdhKDbDvR1P6bOxx7oq3ZrxZkIa/jw
gdmGdB6VT3Wtk5SJECvCjvpkqRCt+RYjZKQuxoXmVnp9sTqiOPKLXAFUviYFVWpvfFaFpSeWE99R
FAXYBn5Vz5cL/K6rALD099LRdOsM7QNvuBBmedLO5D7iOfB4LJvRAdhUutGiDTlf3Y6Dk8rz5iaj
icDvKL0c3AnTNRo1fM5F7+25nsGDNmEHz7zdnD06XP+30ecuxO5cYlKgGIhwggu2UVdirFJMeJUX
C55yfyQe+PB6IVPqfnXAcxoo5u98yUXJgFFyWIriGr9i3a0pDxnyYeBXg9FV36UYajCYvGnKBgGA
JhzqDG9FfrpcH6pbMgfozLvE0wOSIzMFGTKhy75xwA3kimpS8oygYJC2xAm7nmXLLLMvlLpbsORg
yxtSAkq9cddHp8riQdOEM9MT6ntS2IzqwTigXbY4G4DBeVs1oBR2VyOL2oqRdwDnWatyz3U6iUXR
KNsphyLx/ceJSpd/KBno+eXlZWghwlS1a6sdXJpC2x2/pH5b3i3pubWVLlZQl63/AU1eY0GRcM6s
6MCaCBXtRV008SsvXgqH0ccFRTOtgyV3RiLiuU/tpd/XBgF5gQh+L/5A4hD4R5wauQeHW7y26m2I
Uhb5KPUQ3AmHPw/+EgzyTedtUuTE+pGI+XAUda63goy2vT84dLu3tAlDqa/UKhycSnUc7WoOcg7E
f/GrmdLt9MHbMZOmF+NkvEAmdmzYNApolAsc0VmFz3HApy3HZ6Db2lu0dhT6kxtL8q0shHGSPbsi
jk8zV/YZZSFc+uHCWRwwOXLuThLp+R9DRRz7u18VnCO5FXzoW7cwV03+O+iTsBfNYuuLeGbtOKQ5
gQWLixjSq9QAqT0wbYFABemZKO0Q/QNX88yma71d3KyMxpghnNIieGa5sXh4UT/NphFpvOazZuEA
NdzpF+al04mD08eu+RtVv2i9VjPC2psvSEnuy2gRBzD+q1IH9/TYlCQTI8dsDVHNP5c8rcv6PDNJ
WtdGKOl8iUCfiUwPgHPJBdvvQ+3XceNVr7Ph9wCazK1c1yFzre62Q95B7I1SG9CPpv3fDpCDKtbD
8azKxO9FtTxPiYgoOGtCIfdo9YqYAvph0DOgisdg2zApE2mzlZUfsrAzLTeh68b77vrN4Jw+2vId
aB9JcYUrL2lCp7Tgq2InUg6OuD8BB93EAr8jFEmcdLnPUzAC66750oOCI+CAoBNEIMzFnwKb2iER
mz6pSA5xKHxGBwFOvRgXZU23gC0GKzTJcStaS9N8T8CgJcUwQwjFgAJJjobyk3IynqALSZHEnJ7k
lZm0jA5+g+6Dl9r0BpTy0BaWZXjK+E3M8QJyyAlIhq6RrIBCik/uC6tUesHsbxYzwwkBbis76Q6C
R1X3trJX2y6jWsO6iDLnNUxwHRnEQJsX92lvRtUrsl2Asv+HmKeClsfR9o/GRiQq35WIPLiITFKM
4Lh9BYb1k0GxbNgdGR9SfFPA1M3ppxtIgFKB/As0GaRfwKsYp4U+Jitq+Ns/aESF5EXfI7mbC+PH
fbuXaOJt3Q7aN6iBtPAqeN+PueyeUb9zeVYzAXtU8Azc6uJmstNVdctcEvi+MCFlz2r30b3qPyYh
GbWBBtumYWl29tAzta+CLr3jei9PXcy1Gb6LW/hSf/4lDeS2+H9LEIXQCTGJJKKAyQB/g0ucLLO7
J5Iz81+Z+iJs82k5v1jM2ci38lBIQR4IvHZyKITXX2GyggiWFH/8vxqoxxJTjVWvXP16RLRTe0Iy
QkIF27/iFkEj3Rb+h3Dax+4vMUtLSRhReR/Y5uoBbVhyuU6Lzp/pQ/Lv2RjGm6xf0HqQS2MR59lL
Sd0hM1ntrNoHfo1tqki9PUt0OPtUB814CHvQyX12RI4KkZjcdBVPIcH1+cqDrL5e1SHVWhUlZ3Ze
ZDRpCffhqrR06NJYqhGB8fcEBn3mkDQalqK1GwGk2C/N1GA4LdMspttZqTYBmXV+wbP74/BEkr+W
0ak9+2BB7IKN33aP/xOt3QLIos+SVqlD0elBJyPZaG4tljioNsYK3lyeat0jg7RT8RLK0JNWih7e
YjQzasXY4gi1zWzxsQhIEOPqt4RjOjYj3rblhJCT4FQzrWCkmbnkki4sxG1vmF6E1Utf032JZy5N
7A7GIxGyhkT+O4YXE1yA2VLlE7zJbjRf8SBJY/KnHwZ/+EEVzOmzoiLnBmEB//quBPk45r8VoJs3
+wup7ndiUXvAh9oHp1xqvQ7EFPM03GlhjSs0JD37txhtfcg4TEJMUFbb1t1Y6Woe1k5gTsCNyfIp
gd975kfPI4j91Fk/q42XBOG8FAi5TftZszeClDG0DYi2sY6Lqk/lTk7sF8YosAsJQcwjdl1t1Vnj
TeleaJREcxc0BHTlT4ZvRybkUJkb2A4TKYZKa8LM7el6Gd2l+gDirxSefhPKQeIhz8uM4S5rE7Lv
Gw7a5r98BQ2jwzSEfXSODUVSCoo8iqgpcjidhBTbu1lGhfy3ZczOsgzUiSA7VlJa8g+K0IslP1DV
r6KQOcOaBCRm/Nzp8plMzeqYcP12voAm/lqvfq+4As+HLE2LwROYkR6fjkszvgtEbDl8Q54x/R4b
6ty2EYdFjs7NzEAlVooHPz4Satg+fMYevdLN5pMH2JxdAOc0bms/PgPERU4cdnjs1cfFnnYiT+/B
7S5vKXcwoFRfa43Wd2/pLJ05cbaWmaEl338qVFBd8OTPMpmeNQkjt5d6646WqcTYdO15lqAtDFN2
LM4LgVniUj9eG5eADmg2Zl27TGy41Lq5/E/X3JQsrMkLRa18tvyLUf1/dSpiuL0LKMhz24j38Szy
blEUFdA7yz971GvmFjJqVikpl4LvMq3iDhEtV3ZXddfuzU4rB0D3xtVLdUYurI5zfva6eceP711T
LFqnLci/IVVDN/6ufQoIUEMFhebKXAkNjP+cJGeMOuDXq5momgPiox0U3pg8YiwhAxdGxWQGCX55
ESut4bTpTU2gsJmFVQpgyKr3Ldbqj56E8kkDSfLXKRaDm7Jay9NwmTey9J/3XS7Gv8+PlvohThoz
efWlb0nyXr3dlVedWB6zU4OvrpIHrz+TR0QmYCsUUBZc4/mRUbYSKyjg3ECL06/5r/R1xkclo0OU
Ur4EtLgwjGDqMgflVPzUT/SqLV1cKAcz0Q+bUERVFnUy+gkLW1ddxzXocTUyiOKFf0Z6EYsBalny
r8nGlrPZJ4O+qeS0UPKmUN/zhLulurtHnh9VWJrr19ekEILIFMS+PZ2hGYmTPmP7KvNLvBKW7uO0
2eO2XoFQARpYLX2HS4qk6b920MZj4oRzTCRQgqGr2GHcmpDUScLIg25J+mvuUg9mhzRqRpICMZnU
WSM8tXmsJteugZatZexAXgtsBSUkFco3tAZr4xZeGevc/Q6r+qMfaztlkqq4Wn7v3VvzUU+cazwT
SMEsrW+nNQG9iPi1XaTrQK4Bk8JtOPmc5Cl54frFbNQZxMW+eOmewHLgMWOLNtuMe11M4XEuRO7e
owVSz+jWla/Z9nZJ0pnhG1k+CsFn+r5izEBoOEBt5ei7NdxjVyHmIj/XrurnywJ6PlS/NwvcV1qq
wa0/oGngKMiert5oEfYwOAydBrLd3fSongZoMqTI+TBJc88HZ35Iz5/otls6KZRooSgfOPamH6Ir
vWa+ghMZdHTHdqhra4Vb6M5IJCC8t+CSsrz1SXdxjMzOw3qfX1+3Bmz5gA5k+YVxsYUVsNPkHLKl
Q998D6CykP6g67tt8qIhapjiBLZjepJBllKV3+dfe8nfcoU0IksyZZO5A8maMeReE/I/nLcPoLqN
vRv8vVV4IJgVVCq7JsLlBqqnX06+PHr7AR4zT56Dg6KIprcWZ1njRjHbUz79ulQJZtSsmx7+P+P6
m61lH0xd4g2VDXHm0GjTAE+CWUgPYgENOomSCCbbcSPpJq3KjZWXYcZDeULNszM2M++O5N1j0rmo
3cxIqQf/ALFOVFBCN/eNucyla1b+kr0eal83rsw80qYLi9qjZodbbwLsVBXMYoHJX3iKqF26YmIP
skNnm1wZM+YzwOULrpmibPEYHM7hGhD49tMIHckfmKWKXGHkcsgMWnEJBoSsVIWCal5/LcFcv2Jn
DmfC+H0etjaEgbDR8Asvnw9ZOxJUVBQI/7JZsBzhssfV7+loAZfUa144Z85ASmMvonW26iLynlxI
SkIooDJqyj4S++qc5PBdOUsx5PMJuWdMoFWJ0JBAQBUaq8mx7uG/HhAp2zkmX5d8Uvl5vV9I8XBq
mDU7IjvZvECyVc1Rlp7IRYhIJTGzCcHMaOCxc/wBgMqLtunw+hmPG4KPuM7t87zG7u3G3HmBOpQ7
/yFlDSk0Q1mU1fB0fRnO0F77jiJy7ZphX6eBU0lJakjovZuVkfsyUUralU+hrRp5IMf55zaXjT6l
eLy1FQuoLcAiGOdG8xTflmk2dbNZ7SYtmO/EXGDNtRpx7qiobZRK2SI6sUJHDShzJklyLexmp1Nt
pYbp+jQvqRCca3Z3f9n+mrhCBXaE1k9Hf0I/MKvTHxBI4SfZTH1Md8u7r5ONbfouKoahfCayzh98
8B4SfVT/uGsnis/1VFmRO4nqZ+VyMKb0PAFHHmibbFw0hT+YJ1kx3BBVT7DtBJuo7ob4nmrOBxi0
N0Dd+lhtAjLD+m69GUXPguxI9D2O3s5nlVD9LQ2o/mjd/8r/Q1i+JJzvhfqX614UIwpkb0wkediC
rAWQ1/WDEOIrn5zqt1xCZKnzMovQUAWxo4CDPMXDo/CB3Erg2Y1v+t/t+RASQXAU/OCIAKizcguk
vBDL6bi7i/sHEE7CoN403M/wxky/qNPCmClVlSrCGJQfGwlHf5duBQV7rZVMo3B/h3J/vHtUZLjj
ilu0qrJGJFI473lsUwLEzZzwUTaDfkMUaHJn1FRDBku8oh3CGT4nnj2RdU2mqrCJhe/4elHwCS3T
hr/INmnXBN39TAsSlJzQrYo25NpxJmCqUroa8a/sszZKefFkykqPTjFrDlClsfAZBlJi/1XOMxmM
NUsNWQOm1vR+Fqa4FV84u+CrB3OA4ilyrGX5aggdJU2UclTa0cru9zvaKu7n0DJ9+gXeSWiqlBdI
eHo7pHX0/2SEkChJwEHmNqAiyAYgxn4gET0D+MMxsAufAr92l3U/Z7sgNO9rfbyNr5LfqrFnhtO6
QgLEYiB8bNLrjzjDWp4QHcspi4xslNcLlYCWrDIoqHER5AkMJcqsaJgA+T+W7u3Bdh6ESEma6Pjg
NU8FXUuhjVHBfBIL/Q4vBF/7xml7BLi2okvlZY13Q2OmkPJInrquNEupTdQlRNipYK/Yb3SxMI83
qpBI9ch1VoxE4LYCLYXB1IO9G8T/WmS2gorLDbrI8dKkEZrmpHk7rzms7C+/Wson/v3dOjs5x9vR
GWrKnnXO4kUuTv0YwsUVAuatJgpe5hVy5GktOKVGq0Xe6BnCoSvC2mXyJGvtttmpgcfj9KCLL+2z
P1gq03J2mcYRzV37FMlQjGBuDdCViOCt8d2Mc/QTGHbnjdxELAI/cloYlhR59cjzNT0kyH0XLX4W
7jIjYyosuEUFe1GoQj0vy/8g5ofLLBiYY/dprm3aafVBzc/DtYyEhuJEmcFhlzLkGVBfJBWyXD0p
QMCAmRGGjjM/7fNznkskFKTfD4e9obhYc8R16TW8AU+K/zoRd10jsLDU/CLHqUZUsaNOPdVjf7yM
+W0h7zFfygyUHS1O5QfLkD1XsOJpRtP2d+KdCf9goRFxuDLoBO0cXk17aANeIBaQfA1FFrQPwj8u
NmSLCUX2BodhnhNA/xMzbMe++69VRRTJSFmbafiRBOpRAPj9VhDM0j2vb+chC98XfsBlBbCkIMhD
cpZf7DPb5E2sJe224NuWazmILLIXi6sewpbb8vV9feWhbZyT4LEAlZNXTDCnPpHRZVMNkVrB2y6K
2Z8gTFONjFgKFBNGna5Q6aW9Hh/dtwBXXqfPzPGKHuoRiq7vDwgzHYzjQZ/df7DWN/PL+bq6SrSL
sQlAX8xtfv9Tj1hGSkpkwmN87uI6l++BRojbgVAMdSZgjmJbACOq17C0wjgzdD077r02dhLLIfNc
lRK6dz0MKqFOzj+qdbA476lvSV1/ATNLcf5Vf7s2LyYU++vum/FINzjYsTj3NvVBa9fC7w4OAWvL
7lqueQ4M6LL6IvevR8U/YkLbZfsSrZQJApwRDPKQkx/nYBhvnzGITk5zp1e6ZnqpJ5uTWZL4hpRl
GUPGmgtnrlGVFFYjBFua+9RBusKgpfHhmB0LTtvSv6UwZJD0WBNcpa0H4+8095ojnQVAWn5s3Nlt
At/AzS8aOxBQSsU1gsjgCVgvlORHQMPzdOvyVV/x5FYOOqdNvats48KzBBbZWMJ4IcD2qU8oUe+P
U7+Y/Q/lPUb0n+Lf3RsG2wHVHPzfGzroJ4fSr9SdZCUu776lvg3srYhL6g6JNutuv+v/S9PzZcx2
snKPS+hKPQGYXBcD1UEbkID1gpJnegijXLryeY4qOKLagfZidjTMGKOe+9aB3mq9K8+wS2tENNXT
Bkd4VsRHqhnjBu8ULRRnmw7KcsD5AYNMSWk/3GkIDpMULHJtr27QTdlFpKHaoolkGNKc2KMMryUX
iMknv+PZkeNqlXW4DP5IQtSxWhIEJO6xlhKQve3gPdVk47gYRJYuaRHfwXmBcD56Q3mbGPWWaEtI
eRjs0H71u+cLYN8H+xDzyfQ0R5Q8kE6oHHOmcPfgsLG4TUJuG97ZmSZ5jebxKkCEu0Smu3Rg9IiR
svHityv7HWs6paVFjs0h426pRxkKt0pWcFR8qrj7marAT2mKbtg/rVaIgyB7RtBvuunZhqx469bD
rjVVuDflrYa0vva1eBU/DrhBnyeHte+QOLJpKG9CTuyRN48Dv+EjscCMnMKVuqhpS+2AOjUvOcXD
peFWMiBLlePe0xbGOB6+rX1sMIcYC5K/5BlKDVyaqby/JD6m5cABLg0SK3r5zIOXEXvo49M0Bq47
BofzTj2nBUissC6ic3KG3kVf6smT7IkN+7hR6LrYEJ0rUd/EcgbiD76bZifQ+3Gj4Z/DgEZxtclZ
CGHi5dvRZRp/J0jDdXs60GrNOMswMe9eabYKFnqhVNDW3D/11CN9adC/YXyLInVrrS/aVrxLgJB9
uEMUMfhRMaPz7g9PU0IXt7v/FGeNd35V/FMlGUt8eD8Dqd6m+9wXBdau9NyA8CVl7bU1rPWYXt2C
chPaUkfvWii7cM9/WbgzWRlWbja/s74fyhHSStBmHiP7p2k62kNv0NWPfOBFqbIkv9CkWKbDOf0O
boFUNd1lczCJ2lPeB0uxqNitDc8r4W5etO3f7a43JwI3Q8BDWR7oLfbhlLiy4lF4tjEHsuHfyZ25
ZCINzsiK6MY//0WcLFSjgaeCF2MOhQOd4KDphsFXGZoQlQIP6nVv3a00E92MU6nTsZDlN+G7A++T
jgJc8Mlv+rtl7D6GbvN8fjjRiOeaCRZqJ6hSlpgdCxN4IjvjRzJkcrAHhPODBLgrj+bIkwTTnoC/
EVQfDoUyX6qZa8H/njHB2Ni7fMnamhQSpLBi2Bn4vjYbKndQcR5LvbTEvJAk3HYzLVmvirExTSp1
yqVpfHFuRmsn2t9AKTD8Zy16sAWYg8EKQLLz52S9d21Yny2SclYt5cMA/m085pVM7EZoAcbQWbLV
7CTy0kBCULONfD5AQw/7V2hi3LLBxdDXYSvkAPT2MucHn30WRExjz/vdcv1JRup2OFE35Yc0oNRH
gvaksiHV3pQWGP8BT5aN+cGsuhKUZppxkXoFQ/wU+sBapG5N0+ielmJWBNQkqVjCbITLKmY7j2lI
/vGTRiI7sqaPxrRqgyqUGDWgs+k8olGzHg0jY9uurc17tKmHEkvBydyBDH0wx0AFRuu8s2ZINuDV
UpVpX6c8AbwuGb/b/o9jWkGxB+ObliD9WHphcMEWFkXg+2QHN3dR43s0U1Z5sRCbDCIglzOoAX0W
vM+lTe53Pvq2lM3OzfooswrdZUjJjnC+3iEdx8TKBeEl10N37BkrGnB78IcfwLsi1Uc9fR80r3/n
ijEuqhcQUS90lOXrHHbKHi1d6jYa4o5tfZiSytBnngwS+qD9Dkc+eZJ+buwaArJsG5uRpnx/jeRB
6oZP0Lf+HAfsP/3bX90HaAdZNgJZzvL9BDu96A2w/tqrYz4WmxJsGlkenl6OnzK0fMU8ZHUiDesz
W01NL49sUHdkpT3DCVxaIcdMPpHwgNRnFi+M+ME4XCSH/FYo0X4sHppL3cOeLcGhzFHJ+7aJOmQl
GcFE9d2TBHT0PVA4mjVf0/cHdEScc0TktZFAdqPXY4nOYpIM0QjHGnLn3oYVd7Iai4oHQN2ozEFr
bMlq7mNp01HdgjSLgdPm+FNMbt8mmVO0rpE1AwmJTeMvv47vE8YS3JUnBB1dXI1VhFXBPIHNTl/Q
xCmw4ZJvApNUounLnh0v0efjYeRXmSr5qZp4B6SmajcgabVC3jKVA1Imj7oD1uJi80KhAQ6lUW3C
xJPEtbxKTnwlWFgMcTuKRCLiyFRaj7MB7teQkJBQPSECmQiJMHtQEGKZ7kWnUcxoISjz28Iw7Nqy
YkQUqUG4wyp+ZYC2s0jCrd3I5vDSJvNl7epyk3cK77wybAvMhGCCPLO6NtMjYt4S31Gi9FszzdK2
nY7tQ87/dwButx4mt0EOpbTOlCTnp12HbYqoWWiIOL+tkS5TlBbkAvVTg/qHxQcaLNRVoVnoXCB+
MnBvK6BUE+ptrcHmty/vjtrTkEpdF19K3A0jdnjxPq8s5MYfpI2EGDhbhuSDGtOvmsfxjkcflCNv
7M5BRzYu0hXXvNw5ppcsMrHKz8hZ7hMXTlyv8mWF4kgFkcHbI3PnCEKoUWUNAH4GzbgQoa48jDDJ
Fqr0N/p+efry3on22JIYQsvPBezNL6I4JECCOKE6atsNHJlaCK3/CRWcIq07G2nAW2kiJ7nXO5MC
URqV/wD+fPu2Tyuc05S10HwgsHA/3IsWqQD3zUjcEUmjs6imphf0ZwBxUT0w7xsunHchp2JVzFbu
Xznq/CwGRfmBPwvaVJ1VbaCzNFCJDRs2lSIOPo20qe2PsJiu7A1LBGWAL9qFnxP8aoN6De9bz4n3
djGMocVFl0O+k74qJ5BKPhOtZZwQMCrm5noLN2L3OXcD5PodGwVWitosHNOzfFT0+H/wE7YRIekS
gQYZfANiCoOFz5IQQyQE/VNSc01UpFKbO47jOp3QEqaYuym0rwA97krd8nMb39Nx7coVWieUcXym
CrUTKywk7lwdoLNRfAEE4tTG+Cc61A6j2WBhnb7Lsi9N1iuS71l4Oz9+tpararyTyJ+FFHJTgXtz
oIwnIn0b06D6bk7u9U5eQUPZkr+qdx9C8vuE3VUHS4S5Prd8GegvjZKC30xl6o0K1aXBLp0Zq88O
l4BDYpaNR3AV5nzHIdCGea/HuCeuryUXYVkwgyx68m586dPVj4pv+6bst+wjipMYMqPJFRkbMJPp
fJHobIfOfRy9h8lqsPV8bK1vs2CCPez9S3eoQu3MecIK25N+9G33MPYvFasG4RmF9C4l779STHEm
pCdhL938n114m+mFfzjQuBV+5+rRUZVpfeXibG8W83iFhOz0LBSROsXcGQZpZmbGK5rXesbWEQov
jiA7qd/F/LC9NxvX6Ap7RGMA7I/tDqP1CW6js7ebVA79DAZWMARm+eJG2/KrIUZ1Kn4ZSZPaVd+j
9jv7mBvOBdzjs6p1rA3mVRt/ESCf7TfIuWkC/e7A+o+bSDkd2QPFzUvm+Vqj4Q6jdwj60JBOOjK5
B+z9P3B+/VOscKFZ5ecK0TJ1/PGS5nzxbE3KWub7Ef9wjByonFfZifgRAy9cZFd0gO//luJ+jaW1
LSyFnEYkynHPu1gYQiYHwNbd6hGC58HDZIT5fNvkOH9HpYTqmnYg2VhaOjXWNCXO5cmRjMVckh5Z
iZcs4n//lNVPrdo3x1Q0UAIQUzI6wucb6g7X/QJNIYRdppC1ZS3KPZYPCBZvqJJRqDf2/oAZ+6ea
XoVzG2T/Kap2pxxVGGsfawjyPB0HL84jW8MpXmunhvhgskTMUXM/CXCINd50F73BBc6N7XfORRL1
9SBX1EqtqQcWrzat1DXKoXlUvSEkX9yEHCk4Z4b5tTVxgTHmfUC6Z2NmJBxwQPNKfe6umwVIAux/
b/2Ml4NcqSuhl2vsZyPdkOkeq2EOI60NBPTntp+FYEHp/AEK+T2hgX+Vpg4MrDUE1SbAbekpMr+B
DXNeygTFpHUwMJn75tGHi9B/Oaleru81UpFjm/C/yemS+u3gaC1s7qzptHZf/CuZfPyTG86B11Wy
/vPEHHkZcCJ6fhMJP7QXk1SSQY8E6Qrq7IRhc+F+bSxc+SP4PnbzQNStAVuRuUIgU41BHGFNG7j4
7EnIufR+jalUev6q+yxSXmh276kwrQK+KEer3NxhZ2e+yGLiqtihexfEB1jBadJeptRW9+tsiJ7F
xaJGkb4gBRT+HH35JY2gM5kaEkqw6lVKGrwW93ozHGeCInFfbrRQx3SPqUkNvJNlbnJQ0VlDaEql
n9Zap+Qs9U/u5LhiGuLGL5Oyjw48RCoVAHp6VpeKuvx3FtNSnv9ASg/7XV7Wx+gHnaFxZcH5rko1
N6pUQkGwa981lTly85EGSGAGmIA2ycaZt2d0DbsMS/fuFF28W88hVq/EDiA6fS4CHkm0tjZ3xoRl
t81LWtW6tpzQe1z3k9VApo0NdkAiCU1sFaeE71WocdpIQf/EnO5fUkrZGaThfaRBFjKdXLQ8VcV2
56Euxyf6YbqATECFAESfz+PC0OHIxQKVKOpHoilqSZxEK9utYkUD+4+HQH5FWsSwpxCG9CrinUT8
D68xWsYCFlsJaAiEDKvSsoBa2FqUttqanXHnuTmEyQ6t0VVQ1W3XLwTLfxEWerkPyIJ1Jyc5Fr84
pW+gc1g1sIrTRH0Jg43UrC45lDScNPPiP22kn/lQAn8w32mVprxKZVRRK+w+mOl9x7X7wCinp1CV
i3r8/+4zXkKMwD4j9A2Hgry2hpocnTWZLvpmpcs9Q3G+mpEvF9awg2zCSy3tDzcWmt41LRPEDYXD
h0Uu3wFmz3TPs1+AKRzOufzw902N5PDPNabVW/CwxTBV39dn147EfZT1VLBJs7U5inSh9POzhtqK
wIFVBHurgIte+bgYfjYMsvoOqSlprOxaZs0Je2gv39WMxtNl06+OVB2zQ6uZo9kj/15vBziRWZSS
wNFfSiTX2n0xyPpo5WGe5QmwdsZNYEASSz/cNR3De8kwNMboKHC6lmX7Tdb3nLTa39snGERtLGIr
DvnUrhVpK248Skvaf32YPlMrKTSaKSqdLxPqlm5Mt+GJ/Z0h+E6jdspxr+toE7K8k6SPWcwq9Bo2
8mDocHzjmhjcjUhYpdWOzeyRwt6kj/uDI1feFW0SgW+Yp+xOWAi0CuMLtEtnYcf9QjfkvgVzOSgZ
s2dvEt0RYvEBRgoQpxXcoPO/HGZAdjLRX2tNcqCwTUCP/Sa+qhj1rp7j+A9frTjTQYLvBYjmgjJB
Mrk5S5rIMP7fIpC1oQ5FvCfDGW5+Jb2Ddu2nt0LYhqEYlRUKOLIFgc8zmawgh2aoUVIsC+ri42nv
1bMNqtRyx7qrUbIhyXNjRpx254/0PgJFLQCJiD16lPdO5P2mWk7k6A6jglpNvw8vdcO9MZ7xVGji
iVZqk+iWKoOFfDoz52B72C52dxStgAkc8yC3YInW8cPf/SAEnh8v1m0itUjm1X6mSxfSaoKZyyQs
asCUb6L3tp4DZ1HKy4m1e6zvLtCJqLES6L5nyJyOcfkuevJr9dnZzno5jKVqIOX56xbcn8Q8snEL
5k9KGRBO1he9zG4FCnzFYPuzuXdmYk8Tj16+o5e5NISrFzXintnWhkz8SJ3sSzS0lIV/khhnJ0yb
MggZkoCwIDpgq8nPqIlW5/jfi+f5kovD2XtGpo+5xHN2P7tYWMpHVric1E0DAajzAfaAPeIS/STQ
Sue/8oKHfNAqDR3aBH+l0iBKVe7s9X/j2NyJR0147pT7YgfT40mAKMWG5DwuXef3u7q+vjR1IW97
X3l+impuJdMjk9qVh/gECnSM3uGRD/oTCWka2St9thBGqsknBE2ii/3L2oNyR8Tpc9SwbGurDAWo
Jc21Zl5oWmKRi7oxaHYSAMQTWzIUXxRwoQEyoOisXWjH6tXTuV8LjVIy+HMdu0v0o9l+WOqbtWwM
epTnynfyTH8W4XiQd7pqIfbb+W3p0k4HJ1kzDjVxql464fKQA0++1ejsmig3haSUJUESAqQiyMNT
iVp2rT4rnZHD/vE7uLqjDptNgciCrgx9gd+0ZS6qJTNLVt4uyajm2+weu45ATGJZu9blyZOh7pty
zO0ujhlWR7lAUMC5Wy3wcV3W0d7t/DOtDLRMp7eIAKbo0LfveluubrCgRA82IOVO0SYb4woxdp8U
N82DHIODG3QX/+8xXu5rp6ahZHXJ8MgHndLJEAnUqulNA5ttep6wZxEXs2ZrEd9kMBQCwFj26vCJ
ecDCMaC+1zDN9MIQ7wh+jds6niX5PH1KcxO+J+ogDwq9esAb0Q+SbpHcvJXA5Sr5SZqWJB7pQzGM
uXzHl34ILeYkUOsLN6p1K18n4cEgLXhQuO7bKsG6fyUFZ0N4H6UjXgTFoe8UsUHRMcBy00HmZ42B
0cwP1/RtQKPJ7zAHEjhb8F7WNKPUmfM0DzAtQKO0AP05k8bubYP3+63aq2GvLzjLy4RgXtcKV4+c
n5iXVk3kJp9/587c1QCOBohD0wsvA/K7HE6xg3ANUm2B9nqlmLEQQgZE11RlfRwXZuRMoPJHsQ4/
P4xPIBR2v90eL4CcYm0DEfGe9RUFzMj32mYr9zIXN5BJMTniqqBT2/Hnn7QEoYMxDsRjWzmc/rFV
tcRI2pZD4YurwZzVu5D55qlmunlDBcNYPMbgY+FL8cHUCTjvp/Dkkzp1gjEMqbuA16ktpUJ/ecsp
/0lgSXs+Al/u48NG+QzvjBwHTF1XgPqeFfuHlUnjRQvPeu8tVkEg+ziEml7NvwO8GEIbsdT+0kpt
55UPPtziXSJitRxaTGx4oU5v7D9xpVFk5f64UJVHTX9c7HpR6+VRMDF0wD+YHCNYQWfmitJfHmz4
ZpI9yR6x5+kMOLVDpO1ke5gtQBX3fsXV4ezMoMblzqb0njIlSZ05FthDBP5asj+4/ze09pbsjlip
03xc64dbqBmG+S1kX2dutwdeoYSfQ/pW3H+IC9RygAUrKrwlQ7koBCs9AWTd8yY/e5aEYYfJoVM3
WwZYsUzon7OuIdi4p+TQ/KgoGMbd3ibD+qqQhhhbr7QQZ38QLbgwudDkF2phJCnz7KgWGFfRsGa3
zkVU0NcF5I/khdGk4ADShSFfSqZxLpMHF2p4nJSjioC36dsbYNJ2JA4NtbN74SQQrVyEIjjB1SnJ
3chqe6PDionF17w+sqAda5WuHZo/fYn4OkbV3xEpjtVXet9NK8X5qI8Utb5LOnbYUgqHm0sQAq5T
koiSEbGPmWAQezPpmhSoqG1tJVayiDQAif4eDatOeWaTKnMIDMyjyLB94ZFZKvnwNFFj+f4TUgFd
sAdrPIsWx9toCR1WanFeRs2brg+8i3xQf18w4tUquqatoVcyyhuwgc2uNuhxdg3vSX+yKcR4b1B1
BArqdzSF+9uZp553cEQ8rEUB58u55qesh7dJ8aKMNJXyzsFiSREgrPvXLoDpvAjX3kxSiNThoR9z
/Jowg1kMKV16yh3G+EvgFWwQRaReYA0yP6pDpXYjLkzpbd6KwN0Z2UBCcHmYUj5IVLmq1vf4CSWn
w0KDLkiH4wQxrD/nDnHx8C4Q2L5on8kfbI3z9eJ79TRNz8E7l19ePntQozYzRpHnvakQoWdeTP++
w6vWRTJil1mP3SmeM267txgjOpjM7koBY5zPOyPPLjC2fSoVIwGg0W2VqZP6jr56Dcfae42tdlID
tKNhkQGECsXmQoGnkd8Oa0KY21tWrajdk8MienIIEUsZiGuc76q8obVBc1hYP/BegRZmPWyTGFPb
5K/RIwM7JzR+961hZm3+DZSnDI9eLbx7xYuf+CTkKXqwJKlIY+MsGvi4MImLKq6r2qqeVvz0yKE/
wOP6daVFw31wLCC4CRw+V++n/+bxtRpdMNhp6tcyh5MlqY0msngOJQqmv3UYZMoT21cusn1Y16EF
XVpo7RL8Gvzac/8SPeM+xJDbcQBTY9CJkHo+4ClHiWOU5JMXQZsFoKTF6aj8F/dLEvqLgwy1CBB/
M1wwXUqgvFLZjaYVDV/zHkucx/GR7vS2SBP69irFrMCR4gGa61fza3E2sGhnXeBws9/n3M+n1r/c
lL/nzegCpN9o2RuW/yaQL5cSKEjuWvt8JH4xto2htneKe0qgTiJdqZNtH9KJScu3d4yQh8A8DaLk
kuvZiRscRCsmsuC7oZoLLVj9PpS3SicB53xRML4uSpUmQNZRkpaEu6GCHF8fP/tcLx5SV0/L71f2
RBSuSvFiR+HT5ES+ttDeVINb196jT7jqd/mFWIVPP4wFvhOVu0pvORP7bXg43aL61NcZc7EavF6/
mu7IaujufiibWoN/eKDAzM9JNJ90uRRLdxWYw0g3AmccnsDp8whnJm+eMtIoPZQd2RvrCG/2B2rK
Xjj4SQ7KcE8q0Zsgmrpq96/84fMU0q8EaCSk6xFdHIwNGfVhtJ9D7emZPREMzUQvpxqEhDiDnp+j
l3Z7wYzoGxoB3RyQR60BrNNIT3niDyXbYsY2K6Kwd4keHSd0CjgVsHWe9qeGOWwri5dZhu+pbx2E
XnH8I8/gaoNd4E9yRRcAeUaKco/blvHDLkUJ61PUPMV9wOzZiOz74xFiwHia/j6A6SEMCyYKtwgc
OQ4cwITlja+mR8H/sUCjKtXN1nd3FuheOK8iYKgf5CM6yYzi06FqyDZs8/QjnLRHHfMP62VT3m/i
pDSSli0gxjtjCcxaovLXjmtEBVcBAmGAzspAPmaWAjxJP1J0Vb29YbPdcpvuv4HJqprORSb0CYBP
Qp2Pw3Rm3YrJdAE7eLUIhvZd3/0g6K6DwRRhqWNdaHWKLVrOUzMi2g+JKQHH+ls/611AZRkehZwO
pGLJucOK2/LquR+aXgifW10QYNe5wLPDK6mhuiVrJEU9RoOpOXGu/V9xdD7fnDyNe8FzWIsnnYx7
0ucJApHEx5jd3r/v1Rv3QDlIqXfJiG+LyDIJZxTQgZ5nk44ZRESbusvQoaS3PEOqUJTBzSH74swu
HwrcIgo2PQ9dEFO10jMLotC5RdoCqQ9OZsN/U19uNvOW4pBasm1YnYdKeVXCuF2g/QquqzrrMwD5
L5G0WQugOyhM7vOJtNHBDWknAAJffJrzhBi7APR1JBcW6M4bqpZwOaX3KDvF5mkNR4sync0udBHw
B7qWt20SBpNwp4fL6pDnvGfVXs7u3x5iyOBRcm3LzhSTaTIoougIIgTguEG1bai/6SvO1QWl3F0w
lEyL5krIcIwx7zpKuhJtDW4TFI9uKgWLRwreWIVPmPFgMmKVtClkSYflbJoY1QRrSwcbYwfM6rYY
GFjnTmr26r3s0phm1TKWXmj08DRl7dOOD4kyOVWOKpSwwKxHtDlN6/VoknZD7pwk/WyAc9UPdXtz
l82agNYYzDCG30krZes+jbQLQ9/13717lhVjkJlguEVTMMHx90CkI6c70GmFECC+S2XhmNbUcqCK
Zxdyj1OS578+B3KRFefKapX0Yhh+6DfsEBuZqKN643wVsbU0nyPTU34yyqk9gS9aBd2XV60bTSUV
aLo0XN1M5AJOEqCzS+Ukav4FRIQH+thYUmAuSREwOuss01aFGgZdnHhyfsSuN7iiAoFt+X2cOuXF
AkqbFLfQ23LDhz09GplijE+lAKCZsmOZ7nSov7d28632d9/5saSPlS8Oikx5LiFIoCYkCmFptZaf
JT473QXzu2WHV7YbhIolf1mfYoSdYOF+cGQeCvoSDNNQWFLiktKMgwnvvpNURvAGIBc8z/kblzd6
D7/otctJfEUkJ8MYhA+E9NEGMLccHtdmtkHWPuQf4NEvv8MSUWTLz3UOSOmCK4L6wthrj0JbmF4b
QF6jswWiqVbjz0D7SgG1n2F5SoNtl1CozENvtkcw+0Ynk6X/5ZLhWhQUt5MbexUKT23Es4AZ5Dpt
5JhA7PC/jwMeUA2/0sxCi3mzCSWdGpW1CahHQZYnZRaRGSjDXxkeKJpeEyAmZBRSKjJF8rf5cCtq
UgJ5tg4sxsXwm837QB99fOeLU+iSuNnLC85UHCa7/aX8wEgmOIsRNtasuSZMzPxr+TpaO2H0FUJw
iJt97LvbaxUt24iSHq+y6K6N7hZhwDE5sNcgRCZFOgWX2zkdSGjh2cRYS0oVhECaKb4qA/RalPaC
t+HzP9qOOpSebmeDk+EfzKGPcTmGpPERjBI9Qv0fJXy0bBgBgK0AyKH9bF7hY6GJqjgEyCzEtj7K
HpT9YZv9rXBWotidm2WsHQi+zbyeyQz3iWMuUy1YMESS66GDQtsejEs7lzZlB9h4jQmuEI/nAN1V
+gzzq2X9SAp7VgoFKxnCqkhehAuQ/pLmd4E2KVysmKki0EE3Czd9RwJiJ2C6Aw0dyjo9SNX3ogHg
rEWBKzQgT5+t7ElBae71hxAY141GJIJDSO3cLu5I66A68L9P2iObNZ83QAyCVYOt4Yxsa63Uer0d
Nx26R6GwPlbgDJmFReN4VLLoaKt1RZyL00oqR7nQArDTiLxNnH4/cAI5r2Yon7B26FCO+Nz5/+tb
4afWNRSWGbPCMV2XAED18oZFCs7TAdT41lENj1TubKsE75BlMOQW6cWRcP5bRqOvhSjCYnku75Wi
/sWK8Zk1RVWrt8+vPw9zNLn4RDQ44iG7SZsVvjnYeaaCg2IvDrsyHdovO7jSbi/kdL//UPa9v1k2
iiH9gD4OnysG7JzO40GbXu6ls9w2HWiVGab1kFybmuxbzriGIEkiFphwwQNI8GumYTXUgGwBYDlA
24T+WepdRR3CLxucvcGzknowuxVkPaQ/HfPSKdZGJ/vHZP8jeCbpfwQGzflRhfqVVNvLcawQJnYV
lXsJSos1WZrtuWxeTwgd3KqauskMqw45GWgweerXVH+U9nptr3GooI2f4lE5iu2NYenLD0uR1xue
FDEmivJE1+1ur/9AHd7RQQaEzQow25NCTkLSVzW4raBbEfgx1RL6rqoiploEj2ETgDL3ndJBmYrV
mtyhzs1kkwwSwdpk7az9F3yYE+6JxQbVKnmx3rUbn0dIr4mtqPuukxWv782mbR+d3emMAxSS0JXH
Px+hwyrsVOhxMlsNFg6QPG+O6qDeZw0JYrGgrEr2tMuDT3r4BD59O78/wLOfhrbDS63/KEp5NyBz
UEIhArBkdML6pdanK2koHzOSSvvBDhGha1lH/Y3RACuKZ+9mVB290R9pldq4h9ClkWG/2aDviQUK
8DeaPS2mluDH/rPJBgzBh8ETpNjsmZKiyYRVajqET1Udr17Rc0XoGjihSXN/TENPtsNJJXJ71i7b
X6cW3UpSClwO4Fi8rX4W/0W+kJy63JcBixfw0K0uDQL3x21ZLtt6d3RBhqjeXD13Qvbzm6HEb/ik
jPOHeAsC82bnyK6LCTIt3t26SjPmLdBai1KPzRxdf04caJFI83KZG1t5OxHDMVaweENVeD8SDgZn
ZG44gkusfzRC5/ndRTW9WN1AFczCjn6GN3lHLpj5lRx4j77EgiWh3O4nYe26sfkWMeyBLGUXIUrx
IvNdUxD7I4L09NzzvI7NJJvb7G4cY0jWlYu6DkrYcLge4GOpyHOQIdcKxmCgznmeGyD41asvyZ7K
yjSJoSyBjz9LrU97PUU9ouNm5TDdVoRbvqCIc1kyJe58x6nU1tTZfekhp/u3AcCMTUPRKbiOgJg/
afzUC0mt350ri2N5WoSHFLm9vxR62sZp1Ui7s5lsyW71lCZsp+0fN0Xixdxhccd3L2hJcoVQGXct
fyxviVFC7tGsEvoV8WSsVwlegrT/jNw1SMWG8k8YOSQ443yLVS2JIy7nxE53/uLlBSc/XFA5BCJq
LLZmiXh2ioJU6X+2uwVlssLTX/JiMA0lt1FrJcuad4bWmV0WmRJFod4J0bViiIB8ax2UJzTsGcD6
EnbleA0HTrXYHbgWPmkJQqzfE9AMnwRc7qnG6xn18AKAjRfyVgAtt8CUmn3vIEVyE13KGsRWYejl
XWHCHuAYXa1LsJN2ydFm88ZS/I1Ry8A7FbxbAdJCdEi20TdxdZyEvUh3Ux0BQbEPFkuws0gbJ0s2
QcxBP93VF9H/oSDY9cNWZsO3uua3Sm+Nqf2BaIpau7GjbH29Rg+LK8biZ9/dsJv9OofgL3mdMyOV
WsZDy2oKFJamNim7egFvu7rGeMYnJqdCKJMTrOmaBkrbTelfcGJ9wWau2KhT6qbDQvX5jwW2YcyT
JuflIhau1fW2HIde2cQ2wPMI3o7KFd/gYTfv+O9GzrfobciXODA5W92e57jHpkKtlk96fXbKKL1n
jVvEaZdm/ow8DrInW3Y37UdpGYRFJR0ePUXB7Q9T8QOWbpiX+ZRl/Nmw2NXI1RjaDQr+7stmKUag
j0XIga8Noqs2yrNShW6dy0dJ1y4soky6Ta6IArH6Qi5iJJD1xEp4HIcW56o3YQvsKWterJt+rvdD
094F2QfQ65lbw6NJ8oTD9sQ5DHcouAOuQLX0o9fuIEVN3ijw9EB57k2oMF9YYm7fgEQDRWObWdwY
l5ICACET+9U6MiQkrg4R1uOcaLCcAChsiNcSAta2/OnQwG+yywG11Cv2D+d6XX26ekz4asPPJQLs
TCPXM/S3k6TXD+4r40nC9m4CxbaPoBpKC1DbUVYUfFZ5YEFpw2d3F9X05VvhHQbp/vsesKPE6sQG
aoqxGMVihmGu97q8H3j6zU0TRKp616KjhOZkDNQjhtM5Z2+1OrVLtHAvRpFx/n63NznzkRSRjNb7
yPDtx4iHRSGVRcoPBRuP8QL54Ut6Yn0EqW9TcFTqPc4bRJ+xrx6ABvkGeu6OadUrSahDXyJZtBOJ
1HaPyzHxgiG5A/NQMMNlKWyr65fPKbUAkm9MwB1QB4OpnI3kpJSwAAUUgE6FynQSZnCkjby6o+k3
DE1wh4mP2Uz/l0+XZmIakmI6xIbDG0rsir4MYJ0I95rqxdBeb2D8IorqLz/WkWO/njBPswpJBUGB
gWkMtYLX3Yb8/V6YMSPe03MZCWuGl8zN4oWO70Ia8F8cATof31YtaYYzACcgtalPdtVZNhxbDODt
sQWsVfdyYB2TICSzs8NmwTV6BQ817pSvl2OrqnaJ7PGI8xn8lyWHD5Nk9ymRStI0k7BD3+BvGxCn
1Gp05SYWr34YS/TD6FYOXvLwV1qlTFoqpAlQguoIZhE343GX/CLN/zwDdxakao9wf3XRYLy6A7KS
3JtI5aPckFWm9MlY6+N1YMzpxq760EXP1056yonWWwgtyQAJDwdxcOtwcs6aIpWwi+maROdP8fem
s8BGLBxerFk2xU0uHXWSRbdZ7ifuBQSZQUXWLLtfPxpWtx4t+skn4tV2B6kcfVFk6ftgiT3xIzdf
7fSnGM68FuTlnoPa2f9lzI2PqTxLDoSHfPUJILp7SkISUuME59LlRrrR5/Ypx59UTdwCq5aRn9sJ
QbvYrswn77UrqW2Ur5w1i2GhGbnDnX2We+TLPkS8aG32bVoo+tXxe1iMW7vAOiKL+SVkf4MeAMEy
JdWvlVmJLBUmZimfISfdSqywAHHc7aAGNz0Lra7e+RpcsiypJjcqegahWIQIx+d61qHcrepwKnni
Bs/gA7K6quq6SH819vIsCl2jsu+tTWRkPyF35WABQk11phnhAEAGt9tLt0oma53FAi6CQGlCk00C
hFPyBySgTSGs0Jetjl2M5z2NNGGVV9vP/Zd2B3O15q0BKWcBsPk8xHns/3P7aTuMez9+K1+p2AcH
Dj66K7Jx1pVepTIxDi30lduU1DeeHQIgMACXgcAs1m8ePAR7SWemBRc2j38tc0meGaQ+9jMP4OBs
LE7Edng2RFRS2XJB/RHcvrt1hrI1FhAMFl9MGhVtAh1nTSeglJfHfJPA/v53eNnT38qC0lamVXdX
o9/akOpEgsCluOhPs//eXQcyn6Wjvt5dM+X5diaY4EYJgPCitVbgYASXJ0mxJ7C+1AAL5mtX8Coe
b2K7UxFzwM3grd60C/4IlYIbfyEhevRbeQpLb346tquZF3TOoLrtqs1R66cSvplrrx4SWnOBpP0P
1P82QZ6XEKTz/C46W4Y95xTx8J6GpuodHn1KR/to/+rCsQ9YpE/fJInFHaY6MT58VvKpwy2Y+GBN
FoNg5huBKcJcTe1xIMjGYAuVZiJvSe6recwFXpKDdl5s7tOS7Mzd+3OdZ51ZchhHDKZy3LXU7CBy
8CZxaFYdCeNW+RC49D2eZ+j9C4nQsBzWRlnpvlIDk+KTHPyYMtvfiO4wWrhgSVLV8yEObCN6qoJG
Jl4tI/OFKWVPPwoidz/TERcoCqZvuBn5VQIZXHj3xOzmmIUodKkswrhX/4buyMlETgXUUZTaNIpH
XTAdwbXL8x/9LdqE/BCgXwDMbWPFxHoaO/HYvM/1OWfzC6DDn3SozbECLYeD+ujWWPcyf/9wtGHW
1RMRlVnluZqYo05BS24iO+7h7n9j0S8n+WvwGm6nvNLrrV54gqOpXYXiPjxxKSaosgng4swyRCLC
a53UqkXQoczjOIzYtt7bTsA9j0DN5sp0NU5/W+zGa7vRtCW38n388EwXOazUUTGt2qIvHz/YoKYf
uzir/rRl7L8bLoQnqWSapVzMAnanaX1rJXYi999d5qUgUKAfs41IVLusC1GBSLDDD3cuNNfzBwmM
h2E1kf6CumrRk5wpej9x9ps6UMKcGKuRTr5JtJz7kq804x49lAdJVfr67NBKjvlh7Im3uOG33ekK
sOJj6pxt/PlUWaYwZP3XqWenYubpVjDddvbgKq7+DEElCDszWdaMIC/XDSBVAe173NQ6H4RmQkxe
1Pcjbo9brMKpbJpxKpZkB5J/hmJMBrPcvO3ViMyFTjjNxvkTMZHlh01+um3MfqjlEaz1Ec+N6B66
sxl5CwP/hdDG4SbIsInquZsDjHQxslhDcw1mqlEK9oTNyQNydYBykRCxpj7prdDhBRDQyGaCJYif
uJ/cwmgxAhORNxTvdC3lcs7vJpFBlJLc9blzDgplWFBqf+hh5/9jTQn8NUEHgn81ctm6Pdo3bxhf
0/8/ybPIAY9B741bBakHs9BQn1iYUMOR6vmNy//ApiUzSYu3q4TyEQrmj54LSHaCzSpvrwOqnQb8
3N/bMJ3I+estuPA1L+l1KkM56zCAZWUNkJT64J2XehQzX1Qt1Awqfu7Imb1ib0Bnr4Z/bVPlQVha
R7yZuz6iva6gApIiJ3wFhC5XDW6Cqvo4HV3jIERZrLcT9TBl2tJcjRAL68xDkJPu8XjQ+u5GZnr3
TDeNwyQgThWzF4xZjJ85mI1xl29qSWvgeZ5y64fDpWF/Lpgigdoc5D9mMSMI3uYkwH9Okn470Jx9
Y7yBGmSporL5yPWl/hyF5fbldo4LByPOEkxCs1TjEA81z1Mst6thnfdnZhY+IY5GHEtoBSWLluL7
VLn5QgLQmTaO7XnedLoxjGR01YUPD4Sv5uGvdkK0qLW+nDYvAq8s/FYsv04y88ZZyLakK2rLXJ8Q
jLiwiNd31LwD2tAEgPpxHn5LRxl3I6X2Q3y4RNxCSzT8ujkujXICWWC65wXeMD1Bkl0O9L+TzHJc
Q3Zyc4rMMDGSUQLf3rnmvcPPg0QyFoCDqJK0Kd/i1u93I69pVoi5xcMHPbD3+y9Q25V7Ul8xQqSu
Lqgbe8fJEUoVs5OVMJPYI8YlSA9UKv6Y6ztH+whVx83zekhc38eq1ZhwC0NnGfux7AZc+kC1+hai
JqPL5Ltf50c/qS6PADXj053VrnGl92XiZAxL45kSMWSalq6C3N0JUQiaU0q95YPcAUb7HUUydXg6
5BhzlXCr5lwUvZ6nfadM6gdT7DL7eHf/QXDpJHLxjnzqCZaxPuumCDVNKPFMW068xIBRN2peCxED
caer3sbOjqd9A5oXcWu9b7fehVfTRtm6lM6OClnG7mFIomrNY2vsxd9QPLO5al/TfYovfX9dBepq
eNSqy5JLv0tWiG6U+opbtX83DFCxlastTuGF3uo96ipGyG88GikLxGleu8VKUJgu898/08xs46Tl
7H5ln7I8t0ZthfJTz4BqBTxN1TocIDZylTdv0c9fkQHjU7dSpRIHoQhiBoZ2ES2gbNfnf+OMYiaX
3SK7FCcsSZw5abi+vCcvL9JuNGA4fX4RquEMoQ0Xv7lF6wPndYE5Pv3DLcsU73eL1lUxuqUeisZk
xcb/LpkpQvOn9db67lW080DOGaBZ3XIOvL7h7MTskWZgbT3y4+ApR7j1A0dpuNo81sPLETWH3btM
sAXi0h724xxFDL+tkC5X8ne2iglhUCWNLYJbOU2ztaQ9P2DvBqZMr/K/9ergqJsMRSM/7KU3tvlf
lHtz+t/RqhW7HUMmYhYtNzAPg8QHNqv+BhHK4jFuF6N0PkG79dmvM0WCBgTEE0cbTeSSAxY3bjeh
/rqkIpkQ+aZAVo1xrHBNdQvppeS1FvKInmKkuod4rE5EofS4cX3qkDpsItKBQFdZb2aAOwDBhjSH
7egVHeV2MNAazK8zMliSMcF+8/T6JNG7IfDVro4xgpbx4e013VnbjuWK7RBbf3nqHYLOIjzFwDGd
Hx/yxrfJzr7J0xrQCs8Y7NLj+aXUyXKCmVqJxJMByDfi3WcBxHyqinkmJTfSY9MuaACfo+BHZZ45
RWwp1mw26ip1RVqjfFIaS9ONJ2AXsWb/AqGzled9TppTN+j39D8bfvCSD2gKQBYd1eXwHzRqiF2y
y1rVcAy523nSnax7T6e+YI9dYePDfCC6aIYYvnLKN3nftFsjOtkcUTUNAet9DspsLlTwI+0b2c2Y
DGLpXQRQzO2f5CxhgrZXeqs2Qxuc88b1fxSZmCmIkKStqZT4K3pBmmy+I4mYyBrbdk/+jINLLxCv
LWILzxfWijkO7IqRBhvvLrrtlLv0W3rsvDfUn3vcg7L12aX9yTKYJd6qlceYtkKgw9wlLtH+5RfB
EigTHlY7tx1BOqZmDl297VLNffRS9taz2W3/IPiNJDGpYS+GVBt73XXsfINrVu5ChKxODBT/a1MS
JLaET0JgMS3BAreIpStSIVyhXHcPLWZ3EARfD/t7qFGMEqjRBQrwbVY8vWZA/ZM7KAxz5owU8ZId
IljYvYta0Kk/qhumYdB8esbD8YhDQjQ+6Nbqj1BviVf86HDJwdW2gcKZ0qFbUVZarfmilrwhZLU3
4IO+KmFX5vuWWj1kyQSWnJZmkLAmv1Y8ezWC/+8Hy8MrhiLsJqZXGpUgNYOUJ5Ld5XEyaElt9Sxc
7INMey14YMNO9zb6aN4KFtOWMnbP1j3MrhhUgTb6tn3F9eN4V/mVc722bV4gJ68GqQk4NtpnPu2f
BERq420ETl72rr91Y852Mqhgl3kK7yhQ1KWqL+SRH3V6P6jA5LmhvVn5InrI3NeO/VfBVHLDS8TT
sbX6N6hwwpghrM7Gavu1OeRfvvzjMLXJI6TiImUf1zTmE1wXgI49h6Fh/0FJMorh+apHD7scIuqW
Y6Th7zf7VicJ6X4de4IONEcPxA93Hd322RJUtSsE1kij+4eavSuqSjb3fkooMHLeV21aGJ21dEGv
XMCjSn5y7YfrLf/o+UujKRvoED8oj/OAZnjHfAGr1YliqMI577dBXZ2y/53Bx1rJgn8HwgUcpsx5
6UiA6WZjwFCZ4ki58aP05vyqo+8qILxeta+Z7RhmG0tPr1CWIcohtWBJcZfKu9jyav+Rh8rSeRQv
9EgPEe9Y+itiLPaaDJUep6I6u7rOk9Txr+JgSBRTN5dZOGxF/Mmg/ZQtoqJ+30EennC4Cr5BkEbI
k6E6AaMc6BsRuZO1G9evsyKLZUp474t6EHOYVV/K83CIWsMPwYOAwgwQL0SwJvEbbnHEc5xd+hug
WNBUX6u3OdUTJdlPqSpGl+p3KdttNTRovLEULtZ+pP/fIJmiXE7U19WlUVs6sGsA75rG06RoBb+h
kJVFZqFTX39mwrIllyrWZ1Na9wHf59EpUXr5F/ygmUUYd+ZUap8fays4XhYlSx2PNuOaQAsRn8vX
+oVmGpF7uPR+dQPbFF2DmiOtbRNRht/XC7cMYXkdLdae225S9XnH9xiouwP5+V6hNQv6ryFmp+7K
5TNpVu6eB5HhFgAE9EqlOBjTFJ1kXLuLsafBCiX+xQHPqLYXP+9LNy1Vse+TctgMW6jQlu2jzs19
BJlHfgpuQp656FMFZVVA3QmoULXt5zn3msj4a8Qxu4ZMlZI/eAeckU8mt1XaaSgKUvLMr0Ro6rR9
yTYOEh3jD0zRgAUw2GGUBSN7YV3DrEdSAFD/gGON6stn5L7pTJhVJ9pAhhCIceH2ZwBIg93rDs53
vRjIWk/dPs/rsZRsw4n8yKI2f1Usuml4TBczXU6TUIapRz/AkfZP/6JIktfxJjZJr5N7S01QJ6nI
BmCMjl0YhRhB1kgpwmV1HtwRt9DnU8663Yu4S+JjWhLUaRzsV6r/fV40OIyLrgfxyqW4zgbzWjgE
ADlRPCGEGkcuT1Ni3zph/xTyXPgpTGiVJ63QJiUhOv2vJcBAL4ZcHxDLDJlFiUzE8vbu/kLUQ+zU
0B6KU4yk0TYAojCRh9XpjuNZx9OJIQElR6jLB+5ML3bfmURAHF/x+wy32Jf2QXW0kdZkXq8tBPIS
b2p/mj+gLLp/7LPernstJxb6KexRm1VUzgwr8Sz3YHrNpoB7lNeQxdSmeaKZCvRo8m+AAYba+3xi
onmu1olImeD/0QvcL9BJQUwiZSUd5KmGtOM0HQjGMf6kDIzZWI1pSCz4EjV3ECb0mlbmJEvYq5bJ
8ZURzozZKp1Jqe+Ie91SNEV/lUqu9DbE2OmLxwfWw3TcRkBuoQNT5ifYO9wNV0l53Hf2wnP0+6Dz
34iYKqyPQqMsMnCS4dY8eru+80vAVnKfb6wVvMWXpwPbnNcc71zm62O5t18ejJLzg68Widot3sFC
fCxYI5p6q9wHxono9q57Mldt+mKhhIjHNDukgwqPYc2lmqTmAqbfLqLPRpJRPZktkdv8sTmVIFQc
R/Ty5CM2BMDng1gCBSlKmthroTvPTk65CT1kG4fZ57J1HokHKdkHE9/W/+mh2VRmHcqwakaCDxw5
ieZjQk449IRsGg5VdekHw5GpzkxtmkaXw8fcWynnST5wKL19AOnFOUsW26O5TeSBUFtPCCiyqygo
ZpVz3B9TjvUkAbXSgzJkE3wkVrn3mEx1D0+q3VICcTP0Wth7Jc+suMPcrld3vtFe33tBmgB9wRlL
h+3nlQY3HeTQp+D+nA+V5cEn2pGhFsHikx5+CBUWWAhMnTSq8D4p9+2n2vumlCqMSlunxZ7+Ubo1
YfwSvmUY5icvf14gnJvyZihn8GBmmYLPsiINNb38HDPRLeUptitNhD1zOYDq8yElL+//PchftYi5
NckL4ukpyJYCs6RVg8NO/uiykreAUPjxRyau8B9L/AvkU3u6fD0fsJwnMPmZDGpxUO6DAqB3YGEZ
6Plpm5t1ySald/r945XR+E3MsA417oKDS41ZbTz1xJifhy0nU4Z0wuIz+Sqs5c4PVz0Fuj/Toqo/
gpsVGDlDylzVeRLDJtRgj2XsdgRqBBru12Phu/HgUeEYotDzUimadaoVXPrv8iyQC2KO+Fr3cghT
lao9fjt345iWTLGajtoLOFfu9y7Q5hZWAa4oH6qtYeS1R41X5tetHUcq9j/+83N2lwpls/9WykIO
3gakeGGKKniuGm38QnEHd+qlkXw54ij16KrQ+Phbgni0PucK3jSqUiJqGUiYQJPouenpOf6HArww
OULmD0sWqmXdh+q/jnwV2QN01zaci8dHqS9s1OmBhrpx4O17wmOk2Jp4XCJGhgMRN7V3/AxEekAJ
nYzznjFUknDcfBn6fa5oVO0qYO9YpqHOxrK2nF0Zh7yFuwR5aSeEJGlYXc6PTeCgtlPGVnpOMuwV
q9/pDOtswDxkKb10XS6jWANv4sqGPCau5LajHs0k5DRVL9Nb/4bhhDoNZWI8trNl3xImb+M5aRf+
wSWCyygY8I1rY99+5sU48UPjunW1GOMhpXLYCPj3bfA2qob/urkv3Q0pMAlxqaamFMDmxUEwuBza
SYHLzvXX3nwIqHROnJKxn/92NbzZ95RNjP3AMfT1F/1evlDLa9KdesKgmM362dbSq2EZAct9wKJy
6y4DmHBBXKUnMqqb3aCv3tSowefVtNpqFzQpVuZqdAVSPdwh3A7J2GiAar0e09wnv0TnAV7BTmtm
NMw10+KwFXPmQrCNAAua1G7WOQunxrBWJkjQczYFo9a0OVUP/zh1dIbbK2ZV31A4zKaA+BSTO/6O
mgh06BTMBO1Jy55YUrjlCR5/m7LIYIO1PdpnIZKrjzlUkE3gJZ6gbcHK490hMIKQCPEUlYqlKV9V
3UT8btLnUpmwqs2nnQqtsV1oOp2qCepamzj2zCgAb1khTGXJ5lruL1nGDLBY5bI8In4HdedIg+wj
Xyhv4j6gGvA/UnpD7t5/9aHVYgmAjhEE8T6w5lQyPezlkIMYjj7RHbOGMRn/nJS/P0+xvEMjnNu6
IpL0oVLYRYFKymDT5013K0NRNRWkk8N8vywU5Dl4yIr2pT66WuAOykZPJwAoOdsXEVh7ikYBt6Rb
ISmMe29C4yExXMv8k9T78+NpAebb7PnvS1PQ9iKL7gTynYdAdsNhjbJnWk5y19vVocCoJpHsypLk
d02pF4wqWQlKxuP8d2ftpdB+kpZmsSUThYsC93UwuRrGRyZak7uv8/MD0cSwDVEerZaECOVqPIYu
WlFTjUvagRU5OKiOgHArSedcU33BcQtlRH6dUdonrwJRZKK+gT+k8BYxse05LlTuQ117laz2bavx
2dgzY2hVH/AzIV2M+nagzM38wlABcPNIwUFfKNssZBU9Dys1U+H+a+oWFySVCzVgy7PtTf6Yioe+
4pq5rVAXZ3vdoYczdVEvKI4yWTWTX+DE1YeNW62RysNqGu+Tmcxb4eAKKiG1FUReLJ6cHunaR2bo
4GT3Kzf8JbOE050mGln6la7eILKQSGIXcveXQcL8al5bpcWMge6EBijYNOW0z8jCFr5A+onuj4gD
y3ypVui5TxS7ERN46X9Qpneb5Qs0TuAKRMTLBXhUNc4EQJ2kw1GxApMDASqR/812fY5ifu1t6uBF
PoyzKGE6262QngKkQxTEJ19PEwLQd8n4Q9c2GKwpG3/t/wsxszfDcJCr5kV3Hw0HlAzegKOv1/QW
GI3Ft0Y0m6iZfEd+rQmcrYdTkCZo/YMgvmwIDzWvH5P1j44wCq3q5wF1tcYwO1IZ0JyCM+LBASVL
fNtZAZd8bmSPpwxByasolW0LtIkkcIG8JGYfgsl4ylayjeUl11043ijsvFObYRnXZK0Wvg35/mov
kpcbxgg4GBbRmypnyad6KN3OKeytU7mEfizOLzrb9cMFwuu5jbr8xnO5U37/62WclP8Eg12wJjTI
FoO+mFgY/4Q0EDKA3zs4Pjr9lp3+KHDiFAKbsCt9Wx665Ph0OS92qX+USLbG25b7TFU5JQk+cvQq
ltyN1b6kgJ+fpImF5QAcw5mYlQ1Bgfy0nTGPCf78gxuF0E7a7VJFD8ofU3WjoZI+fJt3TN/YOE45
hEVfs+x9UYrlTioY6dSgrTIOp2tNm2fErHYDkCKMm/jWncZzjGeubpA0hNLryktSp3EicivRl7cX
EeGGuQCuSouNmqTqtu6x8Gj5rvn+QDo4qE4k3xWcdq9luBz7I1qmwrWGNuBL5/oGA/gRoHnvfFb+
uWwCU+uWoK/Wf6gi7Dq7POwyK+4kWhPP9Xs9/osuIaSHi/f/G8Vh1+Yme8oHd9jKRTl4+q1rXCpl
jKyUKXTCpDnIkrBvrlHigodu5tyUJwnUyjGUBS56MapXacmMD/D5sVJw/HFz0PtVD310KzFlmO6p
dyB5YVr2GgnBQRbq5/gNue17wA/ohxxzKwvveZ3G2uq6fmaEJI6xi+A/Kl2I/bM9xNi96dhIeNQp
yT9Di9/YYg2pvWf4quPvNxa26rk6w0lh8MFPfc888kWTQvuyFfTCcjsdigcobJTbBfnS+f8/B3EP
bMOkflmESwVk/104Zkei/ZM5ZwIKdfRHhdwRi3TIJlzTdCP8xXaaQ5pM/KeMUrF311FoD1K1jWI3
iOBpERYlxvdHJHObEfXd+Jfqnd3a8O6d3o4h9NT8L9FR4Cc+oBdvwwKsvEizEn8FSamPRiY80Zos
T/4E3xiwDGb/yAivUgsWGp7D8BCjJtw9y4tAebWvfwPX6TP5giCe4BiGc9Hfxt4YwfnbhTdGMGiu
6M7oAYZ1rdoSyoTcqz+edfZOVpmyPFw+YK+6x5Bd3axNvP7Rhw1Le8D9/kmgxoC9BIu1ppiFp1Gb
pXlKjBEVSfV0g1sjE1NGbEiGJYSO8ZcLor3CT5YjzcAIE/rrGGDz/xJqMs+YeSnFVOFOaVIaeDKa
FmM9pjRWNqpoC4WtQfUdrPisI2RcAWpWufXEys7eHuuley3c+FpkCHyEvPq1n3r+/u3RulvdMrRI
gJDMLIr+VogQkFfOqtnnRKlsC5n6/VIyi2ToLp4Slf9xCQkW9nP9yty4ehrRvw3sIWIoM/cp2aaB
pn+yY/fX1BbjWwE3AupqQtV3TUIMHcDDHyfzs6dmuB7736NoLZdDu5XHkNoRtM7RBaQcTBUKzwpm
J6771BSv0Alxni2VQT2MCOL+ruzCayI21OPd9/pMoY3qH+ZZ4stSf2qJ0YYCVUztSuyC49fY5u68
iarj14vwnh6OBoc6sdBDxFhsvrCwitvJvHlTYqAhrp1rjniPwJrHMSNieI9FwqXs2v8N5cl5pxX3
ZGPZuBFIO4JTjtC82+cCKfwu+WkyVyyuGCMv78pk4+lMOvNyTQ8FRtQa/8AOj3/qIxi0jDHcKDCi
2O+VbRn1m2UbW/x6NqMKPbYFM4F2KPvJ+/9kHs/suKsRsb1T0iQ9ZDrgFvtobEwT4CscDBmKHEld
Ozi7ZCOkyibACxS4B2iqDBb73JQK8VeJs36CZpt4QTnethlcPRqWLKxShzsP4Hri/rsL6h8JJql2
lEOQ94dkRaeLdQd5L9LgEax1NTnS5jHhEVJzfvYvOMrRvjb9i5OkPfLJifgf+LaxXSmHJGVIYA0q
KiRbXO7DeSTglO6Ecz1jMqKQulEzDrGmaVIadARKQUPVIRn+xWfxqxKGgfLmC/5PLQ395vbgUUS9
Gr7DptK/Rr7wErpARng5cvmjhDi0MdxpLnyruv1buqzEXhWlHawWX77aMKe51cYsuOyiltxjVDL7
KVGf+4fbYGHtuF1jOckrD60nJs7hae/BC4CxqFgSKahRQiFjaBAy5dRdRnY5hTe3Dw+/1fuN8MoK
jjJdB9oIKvz+8iA2eQnyFqsivuhGYpNqTaNSoj3fU0g9O33tQtCgM7ev6sNIMxCx1i+D3qfsOmK5
tmZeXINjz2fAiLz81AGlk9Tx34fGa9QH15wmKceL6wzIeEsZR0YtfzLBrNkOzTPYeo/UBGk1PO7R
jTFZSijqyuEQa9xXUIS7yh7/K12kWzveZJd1d1FUz67Ib2Gnq/ja3Sk1ijbkZs1zXAAUvIHuM8hQ
a8/zkkD1/IZCnyzAPktPyhTTGi185cfZU/IRskfB0XE5fksICd/KtZodN4w1amRICXQklDHissht
qsHZsLrJAyakXeXbmI4PLMErdauqtjMXmr+b8pwjEYrU1FIJAoQjiYiAkbN6bhKRCLA5d9jEFKW8
C2QNhxn/bqW5FOV1asagCo1H1kJP99V2NIMfyjnjdj8YOBOTdePvnipuULtnBB3N6st5xZXCgLIo
PXsZqRY46uuOSBhPkCzquHBgojTdG8O1tszFsP5UktQa8Wf7EVTWmrM/s7OB2tKuYXt3As6LT090
2TujzvqM2uszPNRlJNnxXAXKjIYOYDLg+d29oVdjs5opt2tnyE5LhgJI1a3gwCXVS1QMsvyFBUCe
tlO/fsyOgtJUROWZVGOuFlAn9+xkVT9qM7ypRaMwHq1ORLaPeBSwIDuad3siHmFEhjozCaH0quZi
0tA60CnXTHrK7Uv8/JymwAtT8Gd72qePn+OZZ1VxrGeVsBSrX5GNCaPWczY2fJ06OpvgXIHvGaqB
OpAwFPKuMQsgC8tiDJRr1dDrfSi4KNmIHWaEdMOQz9r3Jq0dURI18JJUYDiaclhHWfM/t0+2mQAW
MgUoDLz63pqcpS0ZWSbY30Y4WrPzfty6xUFNxdQ9LECTgkj2j6bbbn4mQc+dMT/gb9S5NZE9oRqI
9y45XbRm5ian7aKnku2ugg7dBYs5GYzClzfCZ8rjqaPB0yjnoARcHuhEZvoqjA2larsggYeAZqe+
2DAro8W+Py8BPXqRl28fhId9TidtC/ExMVljz90cOJQOZtkdf4IX0/n9xSc3yoC+YqkmIge1VUvX
NbdiFg5wBLKmklk28zJGkt9vcuMzrpQiP4qm9je4B6ZI8K6AVctBUDLaIT758nat36nSWEBtxiIg
llKI5TBWwVudfqd/GMyx1dzQTxiGBeenm78aw8iD2LTJho7C43oLiGqr4eqZ7TfOVn1GKZD9L8/x
aIMr8SGphos3Ca54NtWycEML/eGgQggfTuzZz6GQImUEYvWDVrfz3acHZ+TZtlBHBsVw9dg6FUyI
pErib2xEp5nWQcszgUB1uPa/TGLfTLkVNnBSm16/fU/GCHui/eEdjttwDSwnszMlBaKleI2YQ+tU
22Ez61jZorOhyz0HXtz2BEW76BuOpjpLPbCH2artgHyNnMp7o+7EBI4YdcQMzPFRBcjN45jI/OJY
C2nuiB9dWUs3rnVBAN2KvAJiCRZ0567o7kt5098dK3LcGDLm95LMf6Q1LwoGV3+IXqOiTgc5bHec
QP6B6xiO3X2JqZEP1LnQRNwmn8l1Ypm1zkx1sGDgEe1Tn4pqN4gU5Os3gpZpTJrE2HLgnIdSWwdJ
ppblLumaH2VYkeFEY2RnkEg4Nl/zLmyDZGh5wmZbgoxovV4LibzSn72ds96/EunVmPvFaNFxBaj/
06miY2XeyR1ZaIAtvgc4EQt6pI1dwCm31tDWnnYkHtZDhd353ta3oC7CVpq8eCDCtPjAKeSmvfDF
yC3mXrigj97NwrPT8fAZ9AHMk/QEIeTTlwEXVPRbLrZco9y7jK4lfyD6LfzusJfPrAfxwyeRIdax
EcH5cN1bFPdJuERrgvMM1/rNA72GKTEdBlS/k3kn0XywZjRvwVKGUN2IfWxF0/bTvHLa66wZ60MK
z7iJXCiK6d+y9tabHema8mY3DK9uzOfVaLxbLtEwWyDUDv8bA1S+JDp1eW5p3r0+Kd0c25O3OlXZ
mjPgUu/k6VHRMdElToGyCXGTmsMfYz6ula8B3fBxYdgrJn8ognfI8wm1Azw9JwHZvaNT3kzoesK7
krx3UnMZItELGuEeo83ogkjeu+cJp4eXN3Lv1DUJMqy+siae8K96Su7427mHBbcFP/8bx/IPBHXf
0MQ3C9wBWzE0FV4hbB3oRs6J5bRDfpR5kYoSWa6Ig8WiYIQJcmmG+pGPOcCNLDj0/kre06Sp84hd
g03XBVnahyghUo+1aGjXRRzGTKc3EZFTavPQ0L06YyKgt9lTcDJQdKwETTnbf49zvGyjIjk1TTxz
sg3sEE5okr5U34pt5i/0mwYZ624AU5XoyuAV5SMjMs0OcLb3ToMvQBvwb9d28m9rrkTaJmk6ov/s
hNjY3QfD23DvLliQcOXw+bRHqHHlXlmXyxRh/Zow1M3hQx+A7tPB2kJy78Fx/+RhabsIZWFfHOeL
8B9zy+alE9KH0mf6u3Yu2z3yLeo9tk2jrET+MHIrgrcwMeSCCMNdS01A4XHFcZu7qgeXNOZFhjMh
yu7NqBwzHFeSp4iXK5g9/y/HhaW41NpERvmlBGWvyn5KcsXg+iKr37g99bTNmbi/8v6y7V2SS555
NXzGPBH/q9XkwnVjSs+rjt5NScsV5g2yoXPLpZLUmdVK6PXU+KsLHvvYJze3VDRQncmjsDHSh/mr
3elyk2McS2WGJ+Qpm5o9j5n0Wd3FV81EaQ2LUv7vnJHW6cPRONA2QPaOaLHvBdeoNaTJUMvJT026
8RLWuE9zFUIfKNYc3jBfbpUgRDRZNYgDeBRl8aUFiJqfl/W2L/dmJp1nR7631sqdcFdwdPQu5IXB
vYj9R5y46lqavB8WVKX5ZN48CH96bg1VL8+s2iMnibbEwIc3ARRUDKRtjSb6XhAme4e/7RKE1Nvs
KPzSyXI4uUeRLn3zRl6kNk1nMl0geb+P+MnYssOaSb4N8vKFGPj+aLA3b/XUwmhYRCb5A6Oc4nMz
3+dknRslPQhwH0EDUzpXSEYUebqMQ59IoeXQR+79444DkhAlbJb9JkObv9ZZS+UXxzN2LRga9TzK
LEQxMVuvUA8BMer63dmko1gH9iIWBJ87sb/OAZJZfy8f35rxy4JhrEphMIBG8OwbfDgoeQgztbX1
FxTaaLY/l46r2+OpVuPfleYY3vsZBA7Nbl1tCdXUx3VsvczomFdat1is9eKQOs6WIze/LCjvnaZS
bPAec6T6JfwqUpZTQ1iPJsAq3y0/VBmnLS6hfjMqMMOq/UGKbBTMvltvhbvj5GIMaexHLDXNWerH
ue57uLcEJmSoTt5YrBnSZ5enPSK+N40onjlW4E9yaXxOlmU9LzBb23SsP/6OsDyHf5kQ7ccCbePy
m043vmBIaigGvMpALJhdVPOuH+UKO2EeTNQB8MyImADjN71VwJ+rFTY1f39dASSjUcWxy6Y08sGy
Wrz2+tdrAci7kMnSmDvBL6n2LuU5GBnBmmL8lVq8Zfr9Bk6Ep4wrtwEpLiK6MSqzKCeLh7PWd6IF
IeWKVngQGXCQsbs/qps/ri9yaKD80PdmtLjO1yk6DqHySnu5nNtJ7r1smU6bt7wnQm2J1pCL5t5W
8HDqfFDHghjFBk+CQXg8O/nzgPK5cvMlWVb+PBmjizIBpWz7eLKq83DRKFYaUQUX2MQiW9boCZky
3VwNpHLZOk0UcuqhM4Jrzn4dHY0lqJXNEgWu+sBL9WZNso8a22Sn85l4aNIX8hXDOxTJ9Lw6kd5R
Et/Xv/NVugBp5UOyXDhEVDNGJwK4j+V9wSpPMqexCPN1CJGutU7ppl2wvOJz0E7FtchdXDeH/GR4
AQiYAgtwa9HrN/LoLnTe2NrSs67b+rrfIf5wAI1Fx9J0SlRE6FpvLB/OapB2rui/SyBh+m2a+//6
RjuVFQhDxm4rZ4JlxzXb22Q0Eogof9Q/BL8w2PR/I1brPutttFiEqH2m0HGHiVFA2uS/aABZQU4M
FwB1EpTWmdGNzIG7ItoQGiXUojSmF7VWyNVXhYQxfXXkUQBAbXMAz9ri48jxsUkzLfU2i+b2jKB9
MBXRXXLPDOXf3GK9sOX613Ax1Gnv3fQU7vn5u41gKRRGqoGkKGZ1Hgy93pwpBBZcaqpeJEX8vSpW
SZK5NMVd22bFwaHQkc5jIWtFufa+Yg7q6zp3dOfgfzmpNk7tD1zQd7SF0+DrUKLkrKXk2k6AFOh+
1It5dLN2iluiygTilb6MXiV2DwhtMm6LAYsp4ZFyTzNp3t1vFawyfQXTIsiyjH4C+xtrI7mrZxRl
wtvWiKM+msWm0KrqZHnUdUkTLVtA/9ybUkarImbiwjq6v5Ar4eXCkuU/3Cv2hsafP/B90I3mOTWg
ajzHoWbARcSc9o7nfWz8UGsgdu4e7YYajkAF152TJ0Cl786SFRg4Ss+Tvp9nfsi0dvmmMV5sx/HH
6xbWrB4feoqeDBxikpfpXcJepvdyiwMGi8e01pv7NB0ICx5vSAKjpubKlhvAUbLz8z8vunnMO7yE
AYYk1MrTDh5J9A9I01PxECaeW+XY1z+oZJx9GtIR5buMnjvYN+hDR/fn8kQ0VMj2T58FzfCh9/ek
4pfVtDSRQoxQcqMMj83dnJkw7ueDD3EFQjWSQeFsM4R4h03TuoN5DUs5KveMbACRFgEo2VXj2N3+
ZR8yKC+YOJZPCRUoGzoWLPNCQBFY74qpbtznAxOlQ4f+uJhrcfaZ9jdflLz1l6wcYooLUEB/ZP1Z
w36I0JQjzzRemq6u08a18+IL6vSqB+U00bGXHtLVUgqNtHu3c0m/kwW5JdjF8GUQkPnnfzhghjKx
1cwGobyKfrQFe3ry4vzZCWqoQ2GPsE6AONsih6uIVyFZ0xbGh70bhct9r+FRZXu5IIc2m1E0xTYg
dP/7zM6DqfOFPoMzAOGoivx0PSpsNq3lwMAbxwfI8QulEsXNyNlE/jn++kWlSJDcQLkZBcF+2NvJ
AHKGQAGuTZi9dB6Q/oM7IsRaRuhhul60mMQj5XQCwjv6vRQJTGpCfyr71/Rigrnq4qgpZ6DIhPiI
TGmZ5l9VvGltd7mmmEyaQtm+Vo4Ar1jFeXdkvqgHok1pETnyWibNU/9q5n+TtCmUI5Bm+KpJ6dxy
l5PFxVq2UMZWf4ixCNbUIYSPGhGp6RwXoP6qedGFZ4+Yhu82C6ufocis78Iu50o1/R/GCVsVVGO4
uFyr7RSIlZeNL9dROVgJWS5WtYj39/60n/pzv5tDyieawEefgVfL+w1wUKzg5Ryhw4byzml5cKzv
YiBoK57NjPVxljM/YjMqHXJpJOH/BFQzvawxtvmLe8UqnAvEiytG4viRC86VjcrAEWY9KDMRizvH
ig64lcRtu8GefkLn+lA2B2N8U3TOUmjA+zzdXAQQcKLdINv3f5MLPmfMCcpJHwF8Af6A0A7aVoCq
6QS9gjgC7l2A8EiPf4dZ5IF4x8eJQA3pMBjS3M/DkvsPKRYuTuW6NDuHxm0HWMR0B99kWKQVMkAf
DSMVWo4T2rRJCaNL1TtimFlpmxxuXWxdTxr0VV258NHs5agHpEH35Wsxa5Q0pqbjCmDyzJPZSmdB
/y8gMuL2pgUPWk8gKse8g0tgQvhk9L/zkxDTKXbPKDbI6NiazXa4o4PFdTz7hN9xO6rdHHcwdPAD
7UeXowC8OKY8+2PhQT/+Ya1UtjZuNF4ngKq8hfPZ8SzDJGGMxe5Nmivr6VI+raUbJV8lGDgB2d16
N0Fb0nFAmhHUXKPr/iCSzrV2OK1B35b9dv5Uff8fhWe1SpV/UUQoBmGnrexaaGl2Zf4Ln88IbxFe
sAiw2tv1MJwhfsL5XJldZYFw7idG8rZuZ4jWMoXyKJsd7CRUMGygz9P/mVHM73V1oWFL5U8rcekN
DdJOEhoLWkW66TX8yGeFHtU/IIUcd8/X4hpJiqfzrOc1btnkcJzvlG4nTbwEjxEasxXvXSgQJQJa
TevbdkzP8fDmSz2l+bS+23xUfTT+MEtY/sxnHQy/BJS21CQrfdg3XnRkHQzmqfp8L0kuqj7o+I9U
ZIJeNNq1bdpA0Uq/nxKvRTsNsY5UnEP/pVfJTtIYMJNruVj4nn0zyo0wptL3cPtvlTbk8CRF1HZB
mfGVxM9E1O1vwmvzGOJtxjGGRd3GMifDu2ab7x+3YpPz4/kyjXgt7qOGV1nX+B+wGEFWZA4WPUpO
70GslYZv+k2EvNh9OB74NV8zHrrJFrMNRO6Tz6TeVTcc1yo36wrkmLLlNzTUol8POoOQsIrcsYv7
eOkCKQFndJZUkJ0RcWN9nCJC0zmgyq5C01TiigwGeDNv5Is6E5usNKcy8oos81HOM2fM3K7H+XIA
EMqxhuo9vCChgb7xUBKaYGe/S3b1QLZaNkYf2g5I84bCkQXuwSmtz/bI+r5j4k0QnWiuQmVurmBV
WRzzD4u6cb7XnvGonBtYSzvv1y5/5JIkcg4ZWuqct1T7fUY4DdJg1nu2KwjUwGfT5lvroUeUf5FH
oHUgQ/qbJC/MNOJVt90qa5ubWl3pMNS6LcHqGsiotLkeNsQ9idsBkl6oe1ry0DZ3Qed6FsqkS2eY
dd9g8fgUP6VvjUiVPLDo7UifKbJfanEB1ScyTU2Bq/YenKwdAGsZTighBtNkjUcrJAvmUA0mW0UK
QI7u8LK8vd2yynTc6UQ1yYRDgqZOJ1g4shXoOtuWkbaVoFuFt9b+PDzEVK4WpCRvzYndg3kw/8pI
ioz+0B3MzBsEmQsukwdKgpQHp2fBHea//GvFCMtFBaXn6o3NejuWk+OQYP0NusBfM+BTRc2f0idF
k4KUUTtYziWOkOMTbv/2r4FEoiY6Osoyg47gO3SQQP/Ctx9X4AfF+qR1Gf7jOIelBQAkCrXAxbDk
vV2mm/iiu3r+MjaFoBrBzLk0GBDBe7xCoZwRzadt5c5+sSNhvSlVdNtDKgtmQF8xrNavHanr4KEe
UVHVYCN8VoNbwrJ+l3ArLT7ZxeEjDxIgZYwTBX9UCBheR2/2hTix+MgJJhHDh7jbyix7/lhkyB4t
0FhvU1wlTLilzznuHaKZhuKYMjYE2cObaz7yu6/1MdtIk9W6WxHu4idcAj+VnCeTrVSU6yY4Xsey
FQfKF1mcgOcIUR/Bo6ZZ+1/pIqnAX1h1rXK23DqTkx35RxS530jwEzsMMYqMtYCgTLgN22FdejKs
cxbLuJNcrQLvhdwDJS+OP9/cBMf1N/LoG3d7iu4VaUJupGWGuuYsBs+bUYcgeJ7Fn8dNNCtI8Avk
6gLB1ev4wjTdq69OaUQ6hBQmtMPEO6uo5zMyRsA823g2aLU3qWVEY5lWocu+E5ABHQ5TCRtVtrNv
+X2ysCL/X2vyDW0wN3eKZijmU4xr9g6j/pudJg8qB9lHUShz5b041qQXTlcOPhCs2aXpq1CUBg4y
Z2U0pA6Ckzm6ujmTeLn+55j/L8oqmduzdiC/PvrX89+m8shrrv23glwLZ8XM2UfHiXkg2aJgpaTs
WqbczwHORmfeSwc8v9wSbMwCJXIlwVmYQJD5RRZ3vLV81nhm0yjzVEakTlw+wzaZ174cSm1z2Ba9
FX+okrzteIiXoniEohL0m6Ku6bC+XPMuM+fU1E38u1Ju9LZNF9/O/jaBHnoJIZO0wFm856mZGGZ5
ENjh0JA23lXPocHwt1Qk3pwNMPh4909xv/WWJjsPuB46znF4W79dgO6S2E1zefix46g2NjpG9low
6lNws9V7FvokjksKOzpInSPuwp/L4APyuO8+utNOj1GgR9f84+u1wWCObSMw65xI+Y09qgZuDJrJ
tOMbjk5ygSaiEYnYgukG/8DecpuybiP+AFR97cSWzmTLurS7S4u8TDMj6e3d+lPJTprwqgq3WbCs
z568nq6G1WPj4KOS18FPPyJSIMK9dbuVnW6ElC4HSOQC+un8Jxjz9FtDy4h006GqjvYDAgvN850D
2iKP6YkwfdJyKGE0ptb7KqqsJhBMMRWwoU/fzOLgX6uf2kTilWXOlLBbsWqlTGwqWTdJYSAaFETE
RyCntd8rdLOmkJ3tIK12cskELc4b6v3sYajvuMb7VYYx7L4N940ChyM5rB3aBp1JxE1z3eORHSkD
EkeM7mwduZuY93fpF+kojeqHtr1B5YzAtEmP9Dgk75rjT2XKdkgwcUowvKTUMub5CTqySlKH5uz+
ow+LjqXv4CXDoqP9G1OYFR/tthARgEF0kOfht1NN3lNuMuSFOxTRYQki7gxJKQNV6hDyU1aYZP1g
9mvfsP7pJfBJ2LYHTWypgApUu6k71v9rr98VIJ3EGvi9oerhBKWWsBUUGIUqXAUdLZVB+L7zr9cP
F6w/zOTu3f8n0UKdYJ9WWFeknVQTFCYw1PR7ZTSG4vmkmPdZzKchaScJSJn1Zx82RpnQ3QTz1zky
puyOma4gtShxzhyVB8MgwhCIdqZKFk0kq+psGjeeQLcGQQPKQeu9ycVn5XrO+G/s766ds8oUU1Mo
wFHMSj6GLIBrpp0K9GVLBLm6N9Qfck9ANGrd8mnJJU5VoIxZl49fPrYpdC3XwWGV97xW8aRMdk6i
MGDj9UTSmwP0urG8clbifkvgp8AOohrjkPsRMYwRGFw8DqICxcVwJb2xeomuz+sm7i2lMr5FnYGn
SU7DL2Vpsh57I5tbZ1BlQUpqzKHN+F9NtD8jycUVn/7HdSbgoRqg+IoTjR35yXZLzrRqu9SEBRmn
ZGvRDthAE1Iljxw8UsfwI74TkUBefqJs1AuYuOHHYu1DV6lG+PcLQ1mKSfO2CNqZlebTNwkLaGWw
CuB+AyD8PEEVE4PajR6sZDGglwsK6sC8YNBKAcIOxZNoqesAi0Zoqur0u059q+q4BzPCQY6JHNSE
CXssk7ZUhCITy+NOpAoaAdXTLY5doeIR1uRcUXcHXEp9sRc5pbzjyuaioyOLCcSmUxhLsGu2RP4r
k85WC9ZBUmS6iQPUNXwMM/V6E0RO3zp0LPoGzkak8ES/RFgnG5OCaMb2zm6LVnKel5yHTSSgHHLN
7aTIae+l9ZHeCvMykKtgA1rizq3vMJNToe8WJIG1/LUoZDwx1aJS81DuLHVmXTmxJ6HM0hVbUao1
T7DkgPqPcurfceJ50sBeToHFIKHpNn3rIRfuT4+uhQ+vD8QCgoHPWiL7H4aoDE+mL0yajMITC/p8
HOl2v4K+NIjfdGDwmPKjYJpNi5xI4pSm3UaDur4ZkgJq9GC+L3Jz1dV2bIOpvEMk7a7ZYN/htYVK
qu3/dIuhluY1MqjI/1pateJJx7cIwRlLOwm+EbRmT5QjTAydIf/Hs7Xz1781/EppVdKNiUvIRPZa
76J6b30Q5WHjdraG6GbHP45sxxUVkzFLjUkxNJn/0fNbpvCVEPMKHPzCtAItetdbiizzfhIgXhSr
qoRh0G1k76ar0wgUfJ/hv+TyJydoXt6yyg1en4ij+w0JT3iGaS3CU698DG6g2MzmmrAi4PpvGk+q
/EVQvjtFz12xIySCyufdLB3el46N95v4diUMKgz//reWQT4NvSDBgBRBiwPqANK/pBBVMJBaTbqB
01EBONjkfaK87S+UisjaJa4hg8mRcgy6YvCoZ13g6YmxNTJQwEiBIkA49XY4YID9xC5LFsmLkjtI
AElyZimkWC1cs+uIg99IfTgRW0XVxoth6p5yQggd247q9qjETUWNP6V0Oxb4a8RXc4oH1KRt+mOE
NXeI3qlagQ2zCNRZF7r5vjKQnKdIIHzk+vS7a1N4I/kwlMN8tt1I9Spj2mrwPkaKDrCsaX3ZVwBR
QZ+jKwu2SKvy/LWX4JdhMicAGwlWnNz2qJzatfADXXKSsABesdF7QJ8JAC3S0noeBIrryIDmDOvJ
komRSVfpKrNkfGtHqqLRWPwWHi0gRET7Dl7o740yuUdKfi7yq4oi9bX+kz1xRf1Cr81cgxu7sLGb
jQ9ZFL5FSGuDcdXbUN8JMx1mtBz/chuhP4qmDKNMfml4i/hvegMY9ILxySzuX4N/f3rsg4AutR7+
nkoXWikL+ZfA7Dzs4awAFUBPR42GEcPEypXwIkyZndjyaSD79ZVCv0iuXX+5qcqQgtJR+x2xPmjd
WIEcuCmN7dE4M86yJQg3NkoNz5VekfZj+DtkOq2Z8Dg0i5vUhWOFKCVKaE9wQ/14Nug9CjDiYVjr
1McNa+O0ZaBaz7NjfapKT0l8bP4FnY6JojnVO7VLRF6aywjjI5ljCexF4x5jritkB/2yVRvQ3m9A
PP6U8IZxxuQh3rwUSBlbLp2Uz0GazXDuWZ5AVCAlqCzSRzlJ/1qaNm7zOh/NIUzUSf4KsQBYjnah
quqmqnVPX9S4D2IftG13YXSmxKkuXHe/3FPJDGC3QxashjJdo/LJSaCJVrvh+VGB6U2Qo/FibKK0
5qxick4oMwSvv+SEB4est7dlRYsZBakBZmP4gfo538Srmu6XjDslTdy3ut+DmDpUqDtP1k3vvD8S
qQ3erwBj1pVB041nKBwBQ9uonhsJ4nWo88xtT0eAgaxQGuk7MF7DX+Yxa7pHY0PhWF4XsH2su5ND
QWES4CWNjMMPYNWhO+thsDD//FQBb1YhI0mHNVMzn/Z/rKbuwBgDY9RYBhK0eAYg32N6FpMq9mVb
ThMxE+2Giqq4CE2e8zu1SRe0r34saQy1e7Ebx6VJG5wWLwk9/m8zYqXozCE86V9uUkoz5XJ4A0k2
mRgjRoTPsns1RAIkmPdBL3QRq9OuYPjzRKDCmPMBPPHaotKZqcwH4pmoNH6K/d1QX9CqDp8JhkyQ
BqcZosWW8eJ84gnB7tfKwc7l0EJV+pzt9A5LugS3Twdf8M9PcQJLuv5AGvwAGbea6qxY+89rQwxO
meLK/wt7V5WrLY447YtJtpYZPEOnRr+QyKi14goV0mBAR7QbxSS32OGSjcT+FoCFeV050nLaiRjr
zoKT3bmpYRo0LeyZhTvcKmBdOVsoVHsvcaNSXeY4f6bDG+IaJRiF4qdCmUt4iRwfOcYx5RLc0mzn
0aAXY57tvt7PXi6XGw8hXUmXxw6m8kV7zZHiqIQnlQy9O69mgo/8LJkqQwTq5Z4D2X+dK/Tuzalq
Du558Yv08OhfcEGmCmquZW97C+7lPVy79Ru5m92VW3/bnIzExTuJfe2EkJYvlY+pgyVNvBA5+UCJ
NIBCTjQeW2hkCmKNEqYDWUNQvfdGUv8HTtzsmonugiaB9LCQ6Q0mc7HCAI3lclOQpbDWEZL11C6d
fVA6pvNWAG6Rp8j/k3YFMJ05//gulSZHJNE2C9KE7w8Tg41BoRiRiEc0cTTXupbSJDUftQ94a5XN
MP/mqdMJmeZda7ibuWPivqCfOVRD/j08lv3qBYPOzEY+32e12JqlsZUgXKk20Z6/sU8WjOEzkgDJ
+6hqvU5SWPANS79nAZehSbvJJLDfqHIx1yLlA0jcfAoFYOlvOyaWk2SNDvalIAYZx/G3e4HDW35g
gD/BEFzRRkk75Z7IgktMoQFd3KH8jgBRDopifllIrCXKnFEd3JthIs5ARpJoUVCjmA7X7wsHgAEg
5mgpjV4z+f8QAZp2+VCQaXf92wPC0XvBJyJjoCFB0ANqDtjH2u2pD/A4/LGVdFJ3Gwg8B8X1t4YI
stY5bOLcvcNHiBCUbjnfdj1YA4vLy7xXPb1oxGiBlN3mZomy0AJLuHF2rCrp3o0b2K52lzLaBH0D
s5u4NUyBIR0+0vHVlIfkiUJ//wFbf+NIfLLLHBo/PW3+0ZqXCsNzzA9boRIB3t5c8hUGX51FviWu
zlDJt2uKOSm1Q/B8ugi+wr5nvgzO0LTvvobBQedzz7NlU5Bfz0vgExb9znpZYQwItADbqlIKrtTq
ujZThCxIezjOvnONBG/pE/Ip5VmsoR+IrCZ5phk0oJBptYjezatDQgQv4DE7mke/wlozhgQzeZAI
JEmTLRUm4/r9ihzIclBWLvBZ7g0Gf89CTT4Z1ZtUI7MlxTR12V041yItSfwfFoQaRM4aMbd+BAAM
WFMA050+AJ6oOPo2/MspSPvhSjB+NAhIHLHjYcV1lCSMLpXPYOjSZgCNUGFgcFqbwdOO7uPuic/J
FMQkEqaR5XFrrErtnLTyZdG97l0QJD6cEK7CeDNFiNnPn8B6IzKai9J3k8f+Jw7g/Aodnj1xqzDR
ka4a/ymzCGO4BvivkbjUxTdDgeXpTDguT5ItJC5S0Jj2DYIsEHIbCmc2W+BbTdKiRMTtD4luFgdM
5Sug3EI1Z6ctE28d6n7FcghEAOIgiL3Mod2GCJw/6XfWMXrZWTU7IhHKT+AZIS9/17hrM+Mm/WHe
vQlPkOc4YnnYhwDkCSCtuEjORGPWbSJUoXdSPQHTXmZjgfEUEI5kdCpKrVpKontYhe8NxFT3OdLY
Qt/ZDcNq0WI8fB0Zg68tuRCmI5Cw9gkH/w20krvjMaeB4vQztXuWc0nM8EmeniGfblmf15B8/TAU
n1CIPm/KNwhOEpHelbzyL1PIOjHG4OvDCkWh/8KkG7wcryYhpATXayTMyPIu5k4DZC0RxCgLE9mB
pgBbS+endPipdjhhA5CvksOvTYXpxGyi6X4pTaUcvJOyNnRoFbGpBdnbZsFrSflQQ3JeNNp8lnqP
NAG4TkB9B743HCS7I7IoZPf+jxs2qeWtgXYYRTzCK5FaJiqaDsB/+hdoGDnKVjX9JCsHMSWzn2NF
0NUPfmGDT4A3uxQm6DcVdbL07RB1KT+kYPk117yU99KwRBCrIjlFIOrtvhjiDvoUtdCancbx1oUQ
HXk9zxqZfLFPGPQK4FlX4BHmc42/3vtxph7bidZyKBOunNaIGHz1bWv2MawZp3YwIShukrC8OKBU
1zxOmLr5FKJrA2C8S1KluSzaLRQMAblekvVP6QfYHfJdVsm6mpHjrA7bSD/ZyDnWnFXyrMzhLwl3
0n2kzDdX4B0K1NcKuAcCcIdGbZWIHmeFMYACREsUKAVyRAzFmAcFg4n3WS8Po0WvCKSote5WZxSh
KCPkn7dV63kTEx1K1RDGJie036CkVNIINwt4e8fn2FbwY4K0f63oD41JFE1G4NF3Vm/xt1Mim4eI
N4fBAVbbOGuvA+kfX+heE7QU1LiXhH2cufofsz7RpAhFkK6zu8MmJ7bbCBK1As/0tuj4JtBN2/wc
3LdS5oFjdFF2tcDPjcqQp5XEJhbZd70j6eNIzkDQYlCy5EWF0+Bc91KSH91TTf3ZP1G6iskLPyZq
LmcFOKcNGOPcZX4SzrJZzsj5qj3aTKrbEd7GiSuC7tRTfLih67CCYm971OE/VZSX3YcMAgTYP5y5
OB/PoZ6DywtAlz2kuJq5aPEDrbVb0XiJ95vS3rwqmy+xmfg8NMNaVMexyrUYzvCHqm6gN8IzJRTK
Og7pufHkUylLIxETl0iVMk0Z6nMNvfcI27x2wBly8x+bj6GR6HKC1RRtmOU2ytCaNowLHtmsLX8I
8+qY2syHGlqTajTalGqwsYaKbdUiz+ZQ4h5j3Ez16IfvLlR7/gxfeRFQQWP3B/3mlYK0E9euxPKA
gdSZoLNqZ5BSzL8RuX2sfr5czoJ0+RLD1YNwd0Y0ZvN+sc0EXwP2iqCCvSnxFTGZknoSayBNKaU8
ugyWsQdx5jxVrPaRhiCLVfHQ/mSGrypcI/qr4NaOEXy0LWHWnYjJqW+UTX0iiS8F0Kvhr89igpFp
A6D/WfZsab9ewBZ5r4WXIpx3N6hlwdzzTQADiEWg8UKglwj+gX3MaP5cxJWVqAviyMsUGus7R7y0
pZC7kmLX5RZUp/x/Ab7ozhqEqKk97AAG749BkAbg9V6bCbGXEtl1yGcd65D6wBM0kjT1rYUVpDFU
3MQEyrFJndQUjDFwhlfr7X4cPJ2gJtMAf4KeKgCNUCHH7XzCpurHMdGnu5GJMTUjl0NhGJAyaBRX
d1up2yoTgjFE38yZFcig67Og+n5pJP5gqedhnKkKk6QxZA4XlwERfxDVwnNlvONWkTHoFuSc8hpG
WOsRkVq5+B3ieHzE9NXoz9dDqK4OaO/ZSb/HGnV/H37St8oGlPaFzJwCIilP65esgdidk4MgCFXs
+6c9/hOtx9/+eGc2Eze9g2hwOUq5u+2Fa+2pOsEz9T5dutQbpT0Jy4TYdhrqfQyzqaHuHdbV3t07
8sE39++E2Wqxj4V6kTS1GqTwhdmCgCdzKn0lBwcv/s3SE3UOYROw1HGj9p/z2dVswacE7z3OpzgS
QVgIheEkcehYfkSe/wYLDR10RAOEhMrDMYPCAeT86otRoDiP5/48CWa/CNuKPYbyfB44qf7FHHkB
nHphHeSWVxNTNGqVkIkiEnb+aQ24kYC1fvMIsPe6TSwwbttGVkZgiueLMkEkvoh9MmQ9FlvKgYeh
jwxZiEgyhgptb600S7b45wp5RdPFKCjqx1lP23UXBrJLdkjGcGBfvd/WRPw8QbTedwR8yr4zd+AC
0VGp4YKZoJRe4ypJK29HaH9CnN3y+JUg2MuEASJxwp1v2/j2kf27msi3DSSdZtnSCBFjL3Cc3ohF
okUOGmFrHr1ttQttq2SKbkkEzwd8ahklwr+v++5758b/AfbizQB32O6bvh4jdpevChMEgxpm71Lf
929Wzb0WLP2N/vvbEhABX+zZT2FljPZ35xhAvHK7mE5wHYJkAgqDZeaWJBVd6wywckwQVg0u0AUY
xJpenDDLwo3cpz9pAQGEOZJaNiD07nLnADUpiSAS/UoUFu1qBr5166OCtiu+8QbwYQMUAhvIUJH7
kW8MRcgZj07eGLVbKF+wx4x2T3pdgygjEITS+nyO/i8Hb6gSAU4jJDSHkwVvuZrbSOByd/m5yuLz
n/EBwrezl5YDL4pVA1X5ZHD235/rvYEvev49k4N4URVbH1IrRjq2GIvwqunfj1asqDP1rE26dxl7
CN2Z1mhqs9IQHcKDUndXIERIHjbEHaEwqv0MFW3FEqaTaB+xQI6I1mghkWp8Efktn561xQpot3qq
6YCm4d0X0g7Wfy6d3aXFWEna04VCvJIAC1ZppK4udB811MFLjY52n/RYQ5qnZWQ31dUzXCv4BgIO
Wx/rNIF48+48LjsAYYeKc/rjJP6uxV4gxfZxfSXmjLZRU5rKZs4/KolVb0Yyb0PfEnNSUqeOwoR6
YFmS8V+34PNezCdECqTFLWIgtpDcm9OChzHhQD0A16GJR22OZlNs2Vk7VNhM/6OlTMhTj+KDjbxG
nzGNm1bkA9ITVWFet4MqEc0TbZ1t0YS7s0zVtBZmDRiX9nintJdUARp5U0gJCRKVMOmlpWEyMTHf
Ot5F5AJEMdKyI/c1ju2LRFsnLznFYVwvZBy+uFPEoipmlGxkYpu4cRvPJYqJ2iyFqOOCsDHWckiB
R9dj2k8yzW6ftVvBL1wWy1z/3/7+NtmMYDmd51iW10aYwnm6kap2nxtoic8bXu8BewbwClrbcmQE
GqpKYPCw/Q1ko/H9yx8io69Neq3PTrOcu1J3Lw4MXRb7at7l0JXspXitMQIarYCv3AMpetFvnAdJ
pQFbCQ2Ed9kZTYxZwJugJITkqLUgF6EcOl/hWtWHfyd8AKa6K2kc7mj/bpcjASMQed3+yYCLSIow
jGLtGpZZDnBr408p8VizAEWSw+KWpChVngy0Sv44n8FDvmSC4BJaPemJHnXLBOKcHH1GGgCFei2e
ucabjYJN9pQJ8PXOl/vDuCfbMUyKs+mkRwaHlc0IrdtIrUSojIJDKDVmDQ+2HeSbC5Gh58lHYrfu
t4WygK06y2sZDZbvRREDH/Fyd+ngbJzNN7Xv5z1/160UYMy/fIqtDqqRHtqlYee0LeH2ku3KfE+z
fMEnb13hcd4dJL1XEm1HpMNLcvSzatUJVibzudSOsDoWaj2kFFjl7ZSsV+z9V4J6oXQ6SJvAFlsg
Bgobl15+tWjzT79nQsaVkEmxC0UlTFmavs2NZRgqwNXH8lQYJWBzpIwxaiLsFAdNvKNEAnIpaeLO
zZw04A00XYLNo/Tiisqjw2qzs0oy7yXHfQB5tIn7EnaMwUfhRxKTDnoYy93jEfXEWSSxDadvFQtD
X5SSwcgFxnGm7q4zpXMUZiHkO83Dz/LBeiB1iT/FSYd8uCFJjqDqmjctjKdmZVRGCUV6rEEZTqnu
bQ60ILnIL9JncKu4lF3EpiXXscSXNlzxoRg3szHQ0Qm3wb1c/OIeKZQjhTkNPrMmg2RgV8XV+/XS
EXGqcGlripjixuV79Cz3DYmXn4S4fR9XlQSHULvlAs5mAFkG6M8sz75aqKLhbknUg3BCH0zdT9K+
lonm86/86ruSS00bsieJH7ynVhjO67HGrP4ugHVpICqu+onu4rwEplkV77rWIRJiEV2RlBdafHrS
d+Wl8TOSABJEqqBj80SKLDLsuxbiSR721PxWKJgPmnIFNikIAHdZ9y9QntlZ5cK59XKAICTodKlu
KSGpa0jFQ4DUayRmngNELg1I5KEs4Og9eSOzgVuy54Gj8nOJTEkJPAlrizw6ozWLhey9y1E03gVR
B4/3bUO/3CFpeoygVHsmL0leS9gZFQy/By9G4oy3sGJJutm1ElusJ6DyIqRUwozNcZIM78G7iFlN
ftVP3jYfKkJssKOzxIvKcpRxXHcI09PuJPZUBbtbFUBp6GOeybSEzmab7+zevUso9JJh4ahPNpqc
u/Irbr/bJkreP0cGEJFuyU9TXtA8ef7zmdP14eBXAaNLKrYJ4uo3+dlCoMZrhBrOEjs8a76t8Oie
0lyKtGePo7SMNkU2wiB9qumo2G0DYvPrt+g6IKbsdqthWmXff6dtzAsMNzXl1QsQYOwt4Rajb5Ol
HjtC1n3FEl6TqP2HzZDuBS65iuDnP6ZHcGxqi5kRsqXrzfMsooQJjILL1GN9YhWUDkSpfNgbPgzc
BdAw91seEXu4ZZE5rA4JPNwu1qluWGjPnzOj6TghjuvMATAoP40yB9ifTPh+JIf/k1nYxpGzU3ee
W7tOblUGYast9O3nj4JEnkplAXbsT61T4sfbMOEFbL7a86K6ovkqvWTzZ2gRFa5X3+b5whjj7MaU
H8o/dqMrq85lfpCd3jbyKlHCcItAvBFHaR9ya0q0B8QN9t4Z3XcYXQi1QQXY2oe3U6W+bh0OIXWn
JdIINaHmqpR5ZoFiD/yEgsBJcb4G/Q1MI2OFLdbJU6tpi0J1AhqccEroILPQM97HA4EzxkMfqX5S
bAjkNjqbvZX/380VpJ+z+yE8/VmSHmXm15puNVlX5M9Ax5Evl/nnmSP7eS7Ygi2t2ww447tvgA8B
ltzJYwyj1hXkxQ64oqhX60QxQdb3ey3O3gG6/d17Z6+qyqfOKcTixEDiUw//WuoLNRVDCNikj83H
8T7MMESmjiKWqIQDKKpdcDh6rCAeMEn0V3AsitUK5ve1xoraOXsSRk61+NIPMgciA8pXfTTvI5aC
55bEj6cbh1t+izuFTleTw8xESm7pvj4quzcBqG/gozWs/UnQGkGnVeXgcvSoSbXnCOgA9kuJgJ8m
2UnoeXd4BaxoyDXjQaJTgkG7NO8Jp2dVklzRzrEQXj91UcFnyF9MCJ1nv1H84DLT3UtMr4DfiRL4
fZCLSdH10tR/BFOZLEUQYg9YNvTb8VvrDqH32Ew3y6y0DcqPMXO2juLbmbyKWmAZpFoo5K651fhA
Rrg/WBO0ecxf+CBav5jZb6bmlmH9pn0ymH1L4Gw0rQw7FFaWPE8qTENQ/a+CETRKPNoiqaVRHbPa
JrTxvFFt4B+hgYsM6JJ7P6BvJi+AFVIuGh0bnI5E++6cAEF9wgEfQlnMXVL6l7PpnV2ySl3bcbDQ
sSFab0+YtTPJr305vyfaYA3VQEEgXZuKIaaXXSZZSK13vxShizIGiRvEpgOpNiV4VQuapgdNPkcE
JVy4eBCsgWtuW9QzJGThTg9QBgr4ksNjjPESUhWHZEabo7miENyJgtDFv/mVJ/nnFgCz2ifH1sIz
rUUdj6pk59WpskBfHetww/aDL9yKDccqTZGc8CYTP0Mn9nVtZu0d3xNsoFXBw3UAurAsiVvWTK6s
wKNxT+N1Z/5+ixgjdeTtn/+07sog321ufPeMz6XQaYj92713m0WDwZz5oh94KWhJvtT9wf2c58Wb
339CMB6fK1vqpt/pHQeg1r7Klvzk6eLi0CFKgy11KY+ku+Aegxc65nsrptCYemLWUWP8qXOSpQej
AraSOeEPW4ryRBS7MDjz2ibXjaN5y+orMEMKoYJSDcykdzZcQO17epTTAfO7cXzlNHsUK9pkRrxZ
PjR7fd+RsWr7CfWJ8RVyCinoS0ELhJprxBb3R52smRgqZg17iYmFdMF7xK0XdAsAXqCQFhJtn4ZY
RrBxoBH7Qo2Bx0FFEbM3kg0/GSSYUihRfAJ/79wHIvbGtOUe4v1peyrTHbHSHJGfPIJODOahDLjd
vtHQVYsdP9egvzZ5RGuvuH3+Sh6SMTqsSCoiHSjN/HdE2vPoo8gRKjZm2zIOCNpKR5Vr59VbR0fK
88aDWD5uWH1mlWr/HqtOtWDelQnICjg8KwEKRxLHf2Icqu/AZv0ZfF8vMNMZch/Fspuf3i8ORAMo
YxnhQJh2VNRBTR0jqbEUHJNfmKIxAmwFv0hHD3LpE8nZhCS25aOH3A6xZ4TyvuD5PaFEG9L3ZLu/
3dUMgXmUzozvS6SDuHMapcphHGG9oU3CPWYIC328dMRRWG8jnyjaC2vPkvfP2ZEhAkT4e7cwE5Qp
YY6Bc5tjiTb/Uzvf7XvTEyHIFm9rf1uFuBthFi6oBbht5doqEmdAPLvjd7+h18PdRhGAR6Jk3Ekj
pOTnpqWuArRFQyAAHsmu+XJLxomBgFDPUEk7BI8D7mjE1FtE+Dcnw5FwnD8KK6PxTUpw55mY2FOy
Gjm40k+sGKtaIheUk2jrZjGRY+JPR13OFlxJFVpwk+Hsn0AyPxO5tFtgdr49qa3curpMsUq819Or
hzZvw/DCcinzcE4Wib4OnjwSS4ysN+ta4SThMV0Xe+I6jFaz0vB0SUYb+1WnOp4YpatCYCu0Ft1f
ytZUeT0FCOhks2mnPSryMYPNDIA7PBPyzIbxsz3wjwD5G4j/8KLLYbJUQu83TEazUN72DmGSkgHz
etXqU4r7dpy16wFKzsTVmRDlDe5I82LeX/PL2kapgwitHUNadbZ1qjZh+92pEGbaX2HUAxkbDmc7
54rAbzhL+u6EYiQ6eA89StR2YzZ8+mYZRVQAbg7KgQYTY+mOzsQe9/JqHUshuMr6rW2XPp284gMv
IAj/dXitxdr8kjtqLy3gAnmOwX5Ta7Os6id6JJWvVnVPDUTBTwQrA5SajlI8Jw3lkxx9TXG4bKKH
7Fe+rENcAa2GvBlv4/uhvVWaKZv6R7bX72ExnQ0cy6zX6uqCXeXD39zFSkgjzm0w0OaBfARV6Uae
AyyHd9KomaNEppDVmq7d+5P3KrjuUL2HW9fwr2gt/4Q0ZWIyq+Put7jgvpX+sOVbrTSItZGC0f5M
yQ0fLE0OTNAfI+j4PfztaM6MECUFwm1VHJbZyBPLc926Xe+oIMB37gu1thpaLqjWi4MhCRLe9lr+
WPYJYXGGm/+46oidUL+UG853D6s9PIkNT+T0VpMrU7V/e2/u1QR5o3qs3tQ9EaB0ZipDB3IQecW+
Uf1evd1iEC3FhJ6Hcv+QAMS5f4Ns4sPS9LyVW460noQF1crTRfk6LQKv8QFBJyyuVqUes+buHEO6
bdXywUKzMivVWgfCgzPzdo2YVkaI2NgDOfyJbJQ/Zjcs9RIid0fWfxcJtLRagE7jI2uKf3DP+6zN
tyh/246uWTZYpmXBu8HjhgJf8EhIVpvarBHF4/iFq8ywSK1SVmcWqtK3qd6SYepagQb71lRx4gUk
zFh6A4DXtvtVnJw/onxqU/v7i/2cSV1I4tBoLrwwi9+ZqknjgVIUj7874n0LbEpZOZfe450omAX8
T0eoW0kNs5Qvgb9yB6Juzp6FFIvWr6oaFnc1xADBtkd6LvpSNiv7prPv0+eD2XOGdc1mymKZ5nU4
sZQDFqFZ3UtK45xHX7nCflUKR5bOqrV3Xdaj3rDJQEGC7mFSrpRnzmWhVNdV1gcKoKuwu+JUqlDT
9lXYa3hYZlAYqLR+qWYxogUEJ6fDCps9Nc6rVXJwyM6GyLeW3pcfvRqWh+LDffWS0SybCfR/pulK
XhRJ5xzMjGooah+wD16VhuoyvLKysVQ6j+/wka1z1OfzBWbaYxXkBohIqr4uxNqhqjpL1GPjt9ui
L3oQgZTiFoZXNULkOp2RAude2fPEwySarfq/JeETm5TxUykGzhulH9X0lsyXqjtP/ehZwEsfL6zu
5HBw0FRUf2PorOt/Wns4UNI+NzplRWeTq7hJRseTl0c3s54iczvG6XPv0Atiy2IN5maxWXG8hf2V
SI/1rLEJZr+IshR0wHG5eLxm1L9s8WAs79d0u+Y1eK7Zmmjg5nKQr62oTwi//zylacblSiUASkZA
ty1NHnqisN83fHRmNEPbMYOnhm97cfhVdTaq0LgrFlVa/x8pUcZV+W3rKqHyBc2V+mHRdfHTZeio
6d9+Iv6OZiwMvBERsPgDUj25tbbUICCQjUBkD8eKHE9QZ3qgh7Ep52+RWoyg6Dj98oo0zVYO/gbL
Jp25rprRIGqQAuNMJL0nelpX9M2HrUyJXyn0jJXmSE+coKAHB0qPqull9250wRTeE7GqUMqiYXpu
Nr3B/hdy/zlEc531JKV+1Ll26BTLwVjqqA59IqIZfHKvuIiacWZ+OyGtrav2IxG9xW7SHdHgE08s
lzazSTLT8tWGX6HT0xJY4laRCMsW0sPPUdPREdyKxkKxqBKkoHer9uqY0CFVKFYTEzKFBNODXcfN
sJZ5eKEKj12sD8V4AbfqefwgOjD96Q+n8cnFAdesZQQ+CnoMvtdtVsKuk2ZCu3gc4Zx0Ic9k5HD8
8Oulc5IrBBwlfPZGW6iNa+P9b1NQ1jp0T6Elj4U/Sj0Bzm38PrLUBXAq09PR/na+sn1XsbB8EkLh
vHQUtab7IYAEGrG9BfsYCoE5Env5G1HJGEt8g5mgNp4Vyz3m2SlzZg5swLXJsDbwkr7vApouRjoy
Y7MzjMLouke5WI5/L+VgzsPbbO6iLOXjE1TUXfTgrGOzxbY9jShv+dzaFpPoIebmVHbNCdZR2IUC
alVMVaAyRd62NEF+krIbq2yfAIDwPSX5PilpGscMMtfiH5WwHZ3Goyb957ol7UNaNrx17NPXhcl2
KZoY1MC5Yn/NEJ1D655Wi0Ffr1GI2BXkBsO1lknTaONfCWAbkz7a1N2C7cH4J+E1HCP6bINZ9zWV
aHehT7CVkwjbLroMnVU8PP1nkR89HE+dQoPFABEtS2VaXSW4HUzYcAUtRiTzd5T3JYmzWzXVKbWT
IT/MQtI5a98GIbtAs91sgAVVlQPdoiT9RxDrOHVnMs0bHKfXKaEJnmXajE63RvO5ADPIZwQMDrRp
IwtZuJisbmdYkLlNwZamjaci62cgDGxh0GMj7KMy12G3LtopncJsJHqq+8YbsBMvGQ6oudXMC7W4
47JwaiA7uciro6QpA2ihkEVr5Bbh2Guda1ms7kKIACkABOW7xHHP0j5hkLOhGk1VEI36MTcPjm6J
/2HuhWp3ND07QuQUiKMrmidZGcrLTMaDtsOv1GLtQSOGBVgCZ5ofwvtx+AVC7uPQqVYrHsaY25bp
j+CsYrASzCEvY/vpDhknxxDNl2DULe0dvYt2qvGDuXGz9lUA+du0Vv+pilTaCpmlFrK7GyKyVz+9
uKvqGRZMFfYuyK86Tg7KG4sLCL/mNut0jYd3o1OOdpb4FSUtI2f0jlLYfxpfBtmEfkgfuaSczXkF
3q/6sPYWGSEg/StMZtgHg2ZQa9HxF9qWjj/odv4fyTI9ttIXQA3wbSWbERxgyBcJQbWcni9KvHxe
iAKlSMqwxWC0e2oZTAkpJrTfc61IrWY7KUQBSr9tF28cnLnR4iccv8EgEdYdZhbZGX6W1ncyzVyL
+yiy2nzJhjTG+FypADW8SgWq+yb7yy2A5TfytqrefTpQk9v4wYKLPbhh4tylbMmy+MpJ/V7B5jVE
9TzizyNvC2pYZZQ27r0R/CxVg/FhqM0urehbra+e32smhl+rb7L7JPtXGE2r3VBK1LPmfX50dsCy
zf73SqkJU958yxx/mLKfaghC1vkRfrMWsx8i6dzW/Mew+Tgq+u4W3UbaE0YRg5Xltgieadpp0M2I
c+1RJzrLDXlH51Mio1FeSHx+dMKNYvvAstjEaEAdk4wqB5cxZhYNvpKHQuBuw7bwWW3YEmfrawti
qy9CQZW0stachZVt4VVv/nBW7e0utTDRxTJuKWVBJkC1roYg7fep5ocf0HV3BpGpJptGiXyl7n6S
kw0PGoA84RmsJR0mjBoV18931k5PR/YT2Dp9IAFfxIPGrE9JzyqC10jc+7ipO6UR4xXfbFgrkSpX
D5LZVFVDQYqqB+963HYQcLYkhITOCzVjzmX1oGDRtecQrqv16tcMG47At1L6BOQT1E3G24QskAnL
Ih1gsoYIpfCWGTzDs6ImFwvLLF6KDKm8vHzDPLmh28vi9U+MskE3aG1wOCZeKN04gA/PJ+dxDi7M
debRlY7PgNEMXuKXbcjqB+VGg7UtIUnQnUvVSUvMGQAqyCoMRBLE7WM8c0duH9lu4/fdDiHCchgX
EGHm6aTbVgNyVdsbFoT/U4nwidknf/OEAAyRoMoy1lIYgCbCnzZ7+dBa9guM/uTRui3QTljOoQtl
fxYihhHPh/6lxvgBESsHPnqrfo250i0YNsH4Pyv358dnjN5vVVXZMnM0TTkgRlYW86NXzEXERjFA
fqzRu+5+LyNtc84UeX0uI3Yh1DlH2dmmD7jxALjpiq+L35i224nzSbqx/CZuX72CwX0vLcBzQIsN
iSxtq8+pxasTdZWhkbIrgYgnQtCaTqSgoZK7PoEKpYsGBQ/RTWFkG8gQJB2//FlpSuWnvunLSawo
t+C1wLYBSzAoT1dSCiWGNNwwYYQSxoPFNwDDU8c5DWI8WnLr7xpfO66jydNPQVyg99HrIrcd+79a
I01GlmI/E/EjsB9V9vKH+/hHu5Ix+iq2YL7U6RqGPAb+DNZQ4fyHlRMtWC0wkfW/PrI34a7pFfHT
/eNpCdDBFCG3+UZN8JAM41Q9ea09YcrO3zpQNiR7+zRGHBeTsCyEmsWIIr+W2XXGNREX6H6bn2E1
xV7S9uTCIdw6GPh+hpVFcb4XUg3CGp71fDljd7OCZjf9gvRUYhXiuU9SCLkF7x+yYj5ODuwvs5ex
GGwDg+rbdm7+I1vSv2yc4ZThAamz7PfsvuVSTMBtY25PdMivSEqBeSbFLOqtXPzjVGwRv0gqmr+P
IJ/x/uOJU5qGyrxj4btD6bbQJnHMv+t+UX1f045hDUpmkb/7yasPdGiO5+KE8xHZiePdtioy7nFj
TGzvjagm1SJfKUFQbJttaGSoW5ap13icN2AWrgZw7eb9bK/NjYyTMXqKcPuQZ+t6avhj6gPIn5ER
CcMUM0YxPZBeYRUmspepVk1wfXGyK8AE633PjICCD0CSqDZakRW+7632X3y9kgB0WxB+g2dnUgi+
Roz8A9w3ibMzc3NNMuFOeH6C1Uxrs5u3R6qNphlpkgyYkfPhla+xkhX+P/9BpcM4/o73I4VCxJUf
jr0LmDa93BR6kIDxXL1o0Px3xPUgaaKRhVkpZ4x7ZrW7sYC2iFR1KQ0fzR+b1bTTSeYfXUtgkhqd
BDX4L0I01QFluUpZ30cQLE4YCdQOO9sEEK4JZZO9Naj4KTdQzC4n7FGJv5tIaFx31SODQjT0SR89
DXjBYcn8tw2OlXpTH/Z5gWVdSjSncF0jMLTnX5Sg8AMxTcTrw6AFipl6jyiWPAYDWERewa4Eg3Tc
JvvJFraKMYAAFqiPdz6tvDr1ETCT0CThYZ5tiypK43RwaoRwftov3C39sHDmm5z3TqaKFEAd2lM9
MMUD3nongj2gfE8kdUJKxWn6yKv7P5sianhoCil//T+lR0c7m7VE9OWV07H/Tr65yIMOUxq40Tth
tBFk1eX7/IkigrlDxVY9sUHGTGlaD49gunw7ZMpRSQpBTI6rM2vE40gJJL3zMbSC0Wse4vHu82bV
/pJekGi7yQy18zriC7Sr1CBw25nhOsgG5w9aPCnUH3DIgnlEsYKb49dbpCQCNt9wBuL9LB2YoJtr
cGD8VdLVGXaOPFu03CWeC5fy7o5L89PjOF/HuDDMgFOCBQdSnSoorpSoKJqeC2bt+G1OWtsY0ReE
iyxcCwh2vtL77JOyJ1A5+M9r3c8Dt5Chb6st10Jy6SIyM9VZBz+siPAZBCEa1An/lWXleUaJpHcv
EheGSiwWqPuX3aeAmoE7zv8AGQN64pT11h3XbJ1UeOdq/MwgDcqd0my3ww+bLbRk7irGykDa9cv/
Bf3mn9NDehLYwN5b1nRcbrZBVNMxGmo49z1OJ2Nf8QkG/DzqEvMqSOy6ILz7+g2n7QQ/bV3H8+O5
yW3i/rnHhD2c9A6RtCch7SxUiJNmGDKWICgz96RqJEYeBRP10r4hJzsA0EJG9VrPWLIN0C8jBzzj
Q8ifHy/tkhdYhjyrMcuVF8Z3/eb/+NP5aSMRbqTEN4nWEPVdeiX3hGpu1F/M8sv6n2bkVkqMp4m4
QOQGSBc7NWW7I/UhGlERwRxKPCAi2gLci+NHszw3Vdx3DODfRNfNQENEujl6YnBYY3EgKm9YVIJQ
1cTeB0Rehd4mYUs8aOm7k8+WiUugY4k/MbW8JtR+Zfc6db967TOYpCKJ5uK4cXDY1arRVf5mfwAS
AQbPr4dY07V6Si/YUplSWOvlr3kEeBIubS4UUE66TvDEj8plZmSgpCh+hdWQ6/CXfFLrrDDYcmAJ
HJxaH9k4tfBEMlKjGE084DSLLujOVMNqnGJZVmkBMAlrXo1eXAZxwDuXerurjxNqlxZtFl5kCgda
40/UbueMjL+9bBGgVmqTAGy3pWPmDZR1BRuz2HVsSs9aqlOKluidVC1r/GGmY+MG3Pn//qApvYdk
3dopmva53nBmXZO5N8Uh20EoWdUwtq8x+nMCg4Glsa9i8uhfIq9SVCV8cfwt8ZoEcjXuK4JBqiVV
+SDi5k/C9TPQt4dsJJJmvheJjAZmdC7QnhHzwfXuSrKMOTsJV0Q46turHRAT9HNTgorB0WYU6bSR
zDzLTSGCUE/svJjR6e41lO6RL1HIuJSSHwhzRlLSLeRYEqm+Pl2XA8SDaG7yMDp2QMZpgWfkUevq
YCYa2oRtQ3HGYD4ci/01k8EFsio5nTzNZIHxe5+4tlrG2iDuhVGHLSg8oDVqpc1Arlao2gE9OXyQ
Ha7vslZS/jTMpR3X3iA86xq9F+anzr9ljBB8unNoasOS/BpZyDUF+QOh2PgQU53AONfgbGPkXT2v
6IXQB7BydZPi3PGrtV+K70XhBwDujA4Hhtr5AmRlF2AeebNWvfWoQwQ6BOMuTuKZswVwt1nIadiz
VI0rUgzkdbt4kG7c2xkXtBwORNn2CWw89+rE7T+hesIr1O5Rka2S+REWjy2ZAip7ZGq+RGbYExJL
dB7YnomdnKrAU1muCfrU/KAW+ciHIwlB2NGFgyueVekn9lg9c3vunE2a4Mvq8WzDCx2NaYzGp4mm
9eXiYp6Prbrs5XYlqDS5mskVvGKErHYPEMDEAfq5WtoshgKAjOn3I5RrnTGsNNVe3lgLbYjui1Ba
TSKXKJGy/4WRLtTRAohFbJTMVz4etXflx+PV/pcfayQufiltp6OEv2GQHsnj4/uiP/WjNyyqwMns
tEmAeSEzwp46NE3r8iMtp9ndJau2/7Ivym9xw6SxULvxWSM295NlI8zGUxuXL0yeWwbl2Q1siSs0
42kE8MSfmipFgm+Tn3VFzlV1jn/tbVgn1coXuvY7rGpXlNssPyrufOGxI68ZxJAjsHV7g6mtPz4/
cLaS780aq5C/PEzIoe4Z+C1e+68WK2e16R+5gugK7A/f8+9NtdBziE9LNNAZDIllNHFZr5oHi1Tp
Z2Zu0IFWM76Wq2LjXkzYsQwIsEPIedcOT84cRTLNTT8IuV2CoiG10HVQazgQg3LXRSETFbxs3CO7
YgXP5KZuaFR0UncV5wnZqAjDM0LPUXntn6xd/1J0T9Gzjtsp9+WaM6jvgIHP4ah4x7n9dKmUC9pV
U8VLtw/v6mHw1Mt+6MN/KRqeYvpEZVZ58/oDbReX05uPuS4cWYZjTufAIrPo0K3Or12IaSaBoTZR
sa1a26GNUJCRiBs6CK9NDp6cJBFxaw3Mt2osqUcj24KXfZ5l6W4d9x6WdnF4PENH2kyAQ/QuIttC
P9Kr+51xTLfeKLCxBbo7eWnUz3wCTHW8XrfIxeD8ZaNOmpigs+CM/UkIpCKDbEzgLmEhPAs6XWum
ESefatpnFmZbiOFKEe+SVZwtSlBxBN1eh0xobIqkbVCYE0VnZXXAIzd8+2mUlySs+pJ96tjKokR8
bcCXNqW2aL8ADETSMdBPH96lP7SlwWRdZylG7Hye15Zwm8P7XI0uxHQiqGWLZplVWGdBRCjDaWDa
8tbduIJF9M+U7MoEsU1dQrNzZ0mDPdPrFrqvFquzNtO3BaRTrMUlF7lnC+B/MzMKjFq20bw03Cq6
5TECEUHxdtkmTOEbbK/T3fbKx8rCHm3Q7MjDj//rRRg8pe3KaOeAVAwEfSxkubJ6SRvI+vGx+vBV
BbQWhijEX2mlSaTW5ZxqhTLEk4mmCqg0hGQTpc4JYJCTsiFMWe08oOp9iSlKstubCuF6wqMiXybu
FjBPYR4RH0jMcjN53ZXLCNO8eO5WKyiEvsfWUfKZBtBlnxaxu0q1OU4vrmwwSCUOvDSZkze9UxaM
kq5mO3KWZQEMkH9PrvrIzWh4niehdwVToEeqDpocgwOx5UE3gnbbH4W1UpkxOl15eOscmbD0JnpN
S5zw3in/FmTUmM4nSmqSl7/bi03aSySecXHmVBCxymx3WCIOHoCC9KK2AB4xJKeAYmsi3dzNzIWz
dQAZNnuC6nlc8nD+ERVsxcZ5uHGLtkf6oGn6lFMKFBOUJziB86CpiRIVgqmWDUmoM0jlCqJ5izTd
ZjPOwpZHfY2vDBwXf9LeBQ02/HWNdCRh9w2LhQkJi3GuywivDYqq9147fdTyXzPmXToUziOJvnrf
eyIAgiCg6NOjIG/yH/T4xKIms2b2/QgzmyvW4sV1hczuZT0Izf+yNFHUphD+vUeMt1vxY6g51Nu1
YpqL2sXTh9bonguoPpFkkwy6VN2l7ojYnczBGJo7SeRZrdBOGjVBsn5mTVAtH1SJqOvJn9Z9/WZY
65AvwcdY0UaOuvwwOcpbuNHwcBzSB+06kJqEoQzpWrnNxNkwRwG9OfA5Qfc1Swx38Vo9vpxR+0fB
BLT0omHYvpZbgRoYpcbsZSZvZQ2n7WWv1tt0WhuSfcouJZbokMDnsRsP96+SsmJhrXEXhgk93dHl
s440eGKvSmzM24xQidvu4cvrTW8UfKRisonOGSy1NsPGlvY5Zq9mbkPORhBb395YfaajjOcCb9aW
GNs16yD6k/DQycB4k/NTEVdlgHPCpj+qkhcjOltMxWHFXIZ0nG1k26viO48Kvsl1oIxBQYXmpkYC
ZQgtX/5/1Yu/GxCJ9f+XuTLKrGSY64JpBjbNDjTPwo+Nl76tAfUiqLfsJg2d/KxT/c6LhqnFguKB
vVirYaMnhy+cSHYlEtvgA8d8W+WgIGCNJ+174sOcuuTMV7qDjHBlERubbbkb0DNLplXgxDW4rQWb
33a6yOnHD6YyW4Q7kp36qeyjpbsn77n5aFYldjCdbSeDtmZ611gv8cEgNQhNPUWhKu/aPPO703vD
8gwg9TxQzdLFfRobpnqsQz/1LMgNeiqJPQXOXxEPxWGyRgQ1LXXlUK2dGKMhdFhwnALKMVWdlTbJ
Y8OSd91dagAyF0JW4UyWI6fn2/+LyDUvF1f9+9CLnjQAwAp5Oaaw6fl0wBau+Hd9dueDAApw+PJZ
dLnwd9hM+xg+BmWqzQ1VhVqzs6lsOlFKvztCeaukqzQGK010SwlDfTQTWlPCcXT+nyk+KopLH6hG
SS+PIUV+FAt4B10e7fEd3GRBexDvYq2ZrbjCLYeInVTo1miC3+yq3KrRtI6u4rRjjH6m2qkUiI7b
/Z2AodrDal/4gQ+mSN/0miAX0fmy2V3xKkojqFUMdHvgW7fGdWp/3muhdSp8C9z3ergfLc9tO7cz
VrsSekB5m++pemOs7xh00cHuWr7iXKQHNGV08LHX/eu9XKkR+q9eZwEbseMCoE1XZ58jrta962x/
UtaZIdMPW5jd3GfhNb/xOumLYQQJFgXoyl4kKKGS3gx3dHgRjzpbUeYS92r7h+kn2OQSOR4Kn05J
/UCV/dQCTOEuutdsvsqDMYcTh4Fgx1jlmJULA24dmRVQUSUjJHNxkNDmSqgaYjjedk8SuZlVuVaz
kaC0eqpXoU6nah+dVSVB5UM3DEygOO7MsksCTpIEPsNaRa/se8fwhCbJZ6gg0fXLxnY58eGlC4nU
Cta7Z9YK2y5Zt8QVqYn6CUfomMLEWAlmLblZap/IjS1X3LFocCGqrzX/5TEIa01MgWXieU/NlmQd
WufmRft+iGXqskGawik4rEtQucpW/vJ2teHrhLPXShKtUsSn4KnV9SAoe2q7eksfdzzBDxQnCbPq
jawJAr7TfDU+/daYs2cl7ZRj0n9NE0Yh2fl4M09u0rqmIdUyQsqDPPo/qTnAVCiiFtyOq4n3FvRm
WLaHMAUQUJ+8yJcV7pX7uRQrjl0MNzNnmrKCYFzlkACgskKnfBLOvfgNLPOROUTIXTyjppzVIvPH
hZ8vsds7/LwlWsA4mezm+fKLf3tiHTfITGrkCG436nyiEaZVLMrCHx/u5mIKnV4vwracUsmfc/3J
Ociiy4N6S+KyuyJQdbUTri7ih+HLCiQ3ye37Ij+RHXCNcHYMEw7CD736z6P/SicVtbVDatiSdwX5
s3rH2c69mKzJx58aM2rBasvrJKamS7tXJi4meGl698LYKc1Y9MPrOHkYSVBXVAVgJB9+y8EBz6uS
5lwjw4aFUXVWTRxi0CUf7f61VSeugXoeBYyLn/c0FsfKeD3v+8kb59ys3qzkLTby81OMA5pXvoZy
py+70SW7Ar8SrTW4c3jJwRMPJrnPpF+ZOUZ0z6U2+45mFH/VKistn9cy7AifxKHPZlDP0gFBkUV0
GZAbaK73R2WqWQVPxpqY0RDXQOUXAtflsku8eVQv0xvPga1G+5t3EtA2YXvTPZ1yttmjrZ8L8xik
dv1GAPHmQJmew7tyqFsNRgcSJz4UMI1c+CEDvFhq6OAuXT51YWRu+AeSKzDaqqwlegaDGjZWUZS7
ATPHE7mNSzYbKOgjUZG5+CjxbvAa5w1XottF/MM3yJ4ngTfc2LCy4uSIzBhOtkXedNi6mZawfFbf
MvKfZohxV79QvacrAKXgsOuXvGtkDGfqNpmJy7r3ZwSDEJPA8bNyfjp6ZvQ27nbxCRtblleiU/d1
OMgmDCB9E8Valm2RAZyaqxVvFIWKb0xPlyhyKORVrBsBWh8l9V7Jn0mY1d9BQ4BCvwV59RSpLRm+
GaHSGyl2Aoo32E8df1t3BWNYGs1HsOQUTZ2UGIM0rqIhct4RCmurBHWREP1krvoQF7L7Q4vwQ2OJ
6vcKoW1t6RuMwlqqRDRaa1oQQ4s153Ks66uNRO7japEpeBW5Xpq/R3MRfBHBlpObMGy8uUQWOkVC
OlK3dHtMhQ2rghMvtGYtfCnb7QqENYTUQpHsoliS5s9MAg2aQ4ZcSrWnjMqJX+FOPu5iztDc8zun
3jSUul4SfqnUaVxnUnmGIr45qutPvfY2BcUMp5Rw14+JOg7RwccqlpSCqUWIVY9OZ8Vg390eEhN2
wbAtrxbuLkasyGq20DET2fav3iGDqBHcCwby7HRdOXZ3I2R+k71XjkcA4BxzkUE8ArhWEKlKZ0zu
fIt8PSVzg8aXmWFM1Vm9HMvgCOXl1mLqthq6e6lmv4+1/kjE0z+hYs4zHMOzARIZDj2A5NMQgjVM
1zU+Uoa76BnhzuESq6AY7cz/R5WRfnS6o2mP42Kz4VEbSrtMqtnEruHDWfpln7hFczyigldpYFtQ
A2ML9f14gyd/wa1ocx8hwicBYWMRIRnIvZZvuybOdGv1h0Zu0ekwHpV+V591I3g8Fxkys5SCwneu
ptADeBQHEDvh2ivRKbd4qWWdNdtL1G0bEbAtIeswWPbKx7DESNMx5Rn0TEh19zmwr0C9KIH/6Ik7
NRWPxLP9oVcucWqD9yt81FBwufwUi4GZ4N66CuvHUEiiq9sEdanEwzrxAdoHrOpKgC6AinMbfIpk
Sm9G5BdJCH9PGd9pJGC68KjtDma3WMsP+IjXj7FjbDoKeHoWH7VEdkpL7RWf08wVicMQu0+vsHPR
WCnlw5oshl+6An5r2ZYXgKVH+JISiUzvMGCzU2emVWSQrt0u7A/O0/vNRwifL4YtAzTmhAKdHLWA
zFMyJtBYnevzyJEJH/Su+4RKAbRKn5TblEEBX2l+k2NjPAjwODfuPJ33Sbr3VeIIyKaZ0Bq+NPcV
TeUNLMfR8F8SxPdH1u4HouxHWrWMgGgjnUYzNZ/PUvov6FtWy8nAD034ycYOQ4AKuytmdj40HJ+e
dZ7qWrdHpioru/h4kt5gMcFiTo2gKVWKmQYRE+KnhlXaXXZJrHK9aeEDGACEXgvNgK8QvPZWw6Dc
Srsf6QxuFz31XcMLkcKULMMGaeC5I4vU5+ilW9eJpUa6KJjypAywp4m4OaqviXZOfryCywSPVIM7
G5lSOQ3ANZv+bMu13iG9cnhL+H2OGMF/1QhUHJY+tAt+Wjlc6UmRVBbOmQZaMc8LGr3x3/wNZnsQ
pSwP3qCq+y+XHFt2Muib+ZCeePzRDPhi+4R/itWo786irQ5mV47oldDRoDJjdKd7UDeZ0LNbbb36
QppQ58QAFw+MfOEqhTPZbR/4T55OBRS4i2ksPjupkiqhIh8wPDBcLfLHFt/O7LmmBD42iq2MLecN
qIEu4ZXDk5+t1jjtqfUzl6TAn5wJjpqy58q81UM4OHt1+aOOZGFRtSaLuUTGSHii4YO8MSU1QsL4
F4ByHMBu9UxaT6CoVClO2VuwJT4ELiwM8I3HFjfXjmEAE1+JoTv6Vnzj4rniA5US8RPLKe2a1h+Z
xvmSXsEbf/zydMBxwzHk5Zr2EDmx7gptU+UcNjst+cAVlYt2rCIzelcWlXdCRvvqsSXfURTIFNUY
sK/YiRrM930cCQ3Un+MrfW+LEqVXM78bDVQ2Qt+w2Cp7W+DBfmKsnoD5CJQTKDTw80e/ZrLLnPtw
KkD6Us83Eq1UO4dXeNjlt2c+VfqxPTdaPaMxNAuundJXVNZLxX76sGlugdxk3g3UG9RcXzKFoDp/
P7HKIMhMLene1HoU5qKAeMiFeuHmZ60wjzrohSVWp1y5qD7lT58KIY6ATbOYk5K0PG5HzR2BAi8z
+ytW026etIMFMaG0BzGfUqpGaScc5Aj8CiViAxCQfWUoh5IQAVqGLFAk9GHyb8KKcUas9O5NFjkN
OlrlOYG10H/h49SEesZWIDxYHkcZaYot1xYPTLT7w50dU+zPD9Et5VG/DtXkovFf7PRi9VaK/tTB
cWOEYAehRzVFmeoisZJ0yjilcq7nhUjGYzfmusouG2CwIo3Or1uG2boRuL3X11CE/a2IfnRZZ+uP
+bYIgCPaDyclioYz4JMCuUD7RJJT4sXD00F7kAPchy7qK+OKnNXTo+a+x5z+BHn3y925f96fEshX
03ROtp9AxH8fKui2yGvAaiy4AiPLP9kWmuDh81gRL3QjhCVEd6VuViCElqNO3v3pjMM9pUV6pwU2
L+mROn8zCBCmXa2fnJi9cV9SNLcKILoJrehJr905O2jrlYK3SuawRv4yWElFyoiumqHTd9jFs+Xd
L+oUGGAb0N5Zm1oKPJdE1cLu55JmbTbkPfkQ+FfCBRITXzncNc2dYruSFwf0+O2T85bF7uYustxS
M6O2RBHct9E24k0PIfjwkOdMsjoCSLeL4uRHuJ5JD18b/Hn7VLYlJkkXZUMfSaVVkKAcAleEiIRq
GzrLC1KO3sQ+xZlT1vCKgq960sF1ugn8fVe1g0nfkBdQZQ+U/BvpUFF7OakrwfnH1oWjfvoK/rNe
swF9dHC63uxVMh6HbzHW8xrCDmY54/jTiCsbHA97ipnJIAlnAhwtqmIxKLM/+Cq8PUvq7txRWJ8n
jEUaelZmaBg2oxWHtbM/f05ZQ7GL3ne3LRgcC74fHEdEUQUGQ6xTq695QBvLSzygKThkuQGDP7kQ
V7Yj+QxMtCZouJKRKQJKO+Byx27HhDHEmf4q4UaFQD6FBnot8sWwtx8wPlwHbGVcJfquALScvhsv
oZIFZyEdvFKVnNgi1lzbKr+IsqA/t5dSvb96G5b30rNeYm5c+MFABWkmh2+KfMgmRbOQhoPc3lnq
X9lalPiPMuTZ+1KAL3VC9TAU9l+pxa+/ATTeotLbb+C1a8Y79qYGZw+mOf1rKil5bqYZSNx/eewR
5yhe0j7J2h4WXWfolBCPxe8r12iJetiixOebuW5ELji1UG8keW3hFT/vilkYovvAl/8D2mp16u20
cIOHdSeTh7I1GhQMgk/eeQJ/eST5yZKu6ofQangEv72D9zfy53bAwhALE8j2w+9YuPIDbpuHXCMa
Oqu3tRCmlC2RKMkyTiY4Tk5T2CkXJsVY0q4P7zwJl72skoPDrSKwxlMKW56jbkW53P14iuAoZ3hA
ds1em97lcBzYA9GimhMT02yeD4hixK/idDYF5xAjdgEM3Bw9l6VVi88KspTmu6ImHER3Z9PLvJg+
Yq7ddLL2yBMVvHuKysjenUxRihozePPa/8eTHzQv2kGkrZudRRYEfu2ntm6Z+SLpbob+u/+H7Dpo
xBZE47kDhaap1YGM5+rmzqgroAFM9m7ZFd95wQD0E7eqvZQGijy1LB5aXZsTZnLz8oDLC2j6cKuo
obWOoD3HEn1RCfwydpdNl2yEjhEdI+cfKH82u+HaDXxdO8P7bUs1HMaxmVKXbtKqp3PLgH0FU/7z
h0fy+38CFWP9nX2WP/zzDmXFfHIyfbSDpqqmxH0DQRQ3W+vIomS2ZmhtTvNfp3oRVxC42l5TTYi8
EkzMAhge4SwRmNy9bOrWRgpdpT05DL56kewDTwdeowGKrQagZawwPiYEzA9ADiemT+MQr3dsxxs3
hQIfrKVR4QktNjGoyWRIjF8JfLKIwf8ciUUFxuaQMOlxgdbKIqdMCGEW2FrjEg5c7k/vVXJyHpTD
2sZWw0ZUalhXgbnQhpJy5trEItYQYA2TXnZsAUs12KWL4jVHqr1sD9SG3k7kDsOmrBuMHHEc99IS
QXwhTEhMflEmTqUfieTNXjsQivLW+ZPp/xPAshbLxE2SwUA0blXOyFuy0mEz7ZSkkHGqCmWa9Hsg
bLxhRp7i0WKWijj9FStHG4bJSLSmyJBnnxWjarwC9FkF4TICi9TnDc0q3NReLmtfL67KPCKIXbyG
5K8S5o/WRTqEUr84tV29HIXFifqZeSqZHwVwMs/F+YoDeDRcv8OQHNMBEoecL/pIbUGkFlN4lgqB
tnB45CaOO+Cxjj0TvFYIFrIDBCvO3Pe8xEnbthQVUCYCS3Lzm1fIEvJSs1QwFOBbetFoLEv0zd9M
rqOno1UUeG7Sn7RAKK4NFZnVAx3CVnC2egB8rueG7qs3QS9vNUWztzNeGr4plnOB1AeWO/96YPSu
7MwIsU1XdArW0xKGioFj38AC/tygavQrKwksezjjHHh1Msm2J0/R6kymJhxJZ1JhAKcYydE1xpWI
0hG+9gqFJw4H6rVPpfqmmb+9FrrUUzjTQ42K1vcMJBYsdLZVx7OMhWdgr2XiU3SqWbOFTvsaq4Fk
lZsgS+Lz553d5F83xPXBN7r+UulkWvYVjItilD7T2v6gSWClCkQbGhGAdY6anS7TymJ1uwX4FUOC
JOaor04ZDtdm1omRpAmOvVtVYMCJLocvSyfRfGXWJIP94ybxkzXKfXmEdfk/t0/VK/DUQuUVsWLo
xf4y+P9Z10sEhkfjn/qFhadVOlS5COi6xSmqyXiQBFh6D3fxfUFYD52C04nN0eNU6j9uNlDIFFpF
fjdCEsXCbvkhVSB0UxjocD9ScdNLmRVPx7ZtivNDT4wrKnIjrOqWgOlxeugL/XB+kdwSwFJVW6iG
DGR+eebo24SVNZzLv8GZ66dsCE5JxgAWT3eUDKgKUydfijQI62vB3vAsA2+RXA9P4cXa05R+7m9J
pKWsHfobK4UUbNgeKCFzeF5B9pLktFwsegC4fzKVwpb5pYhMiESwtN8CQVmzY4JdBCwKNLkPSrY0
+/gfTvqbtpJevPrUrgnja+9XtKKMFyFX2b53yZU7eOc7DMcEsUQL7VgYd/cuD3bwdFnv2kEQTZma
WsHZ9zdErJZzGIn9sBLViUBL1gAOZNibODXPCIZE2/NsnIcTS3g8hYSNBOnbn2aiUEhHFFrgkckm
9fMAJF4MsCIRRqqn7fy49Cm1TsFvE7hGKX/Vlc41bexHMcxsQpB7M+0gAwtlllIs93wIZ43vlxwv
O96DxmOs0oL+RFqYNehezq+FkVkW9mztOFPLG83NfvQ/1Wk/zNRSH8BfeVoI8yKHBnJo2MflE13Z
yoFM2CNYY/sd2tgWtuilIXfEO/fJ70eZWxR8H1OAKKPM3of6SL0euSgbShqLwapTNyUISQM61yq8
wlwng7E9ky+1ouJydQZhz9lX22CLEZGp7rJdAzV2TLvndTBBM0ziJxAfacxOeH4+HDrwxq66rwfb
brQcefLGkggljIirmuoOWy49gADvFubrvHrFKp3B9Mi8yJORfTkslli/dLWkOTw/y3dhLmdfaKRn
8njuFghKE1eT5vKM/566Yftoc9m+bpX4inCib4yPiv0xbLN0SBUwF7gDAKdTk6fqVqzDjVwohKy7
gE9jVNhieRuBhy1KmtgOrgmT1s2tH20Lv/lBEPa+KJ2hof3ZPs7wyKHEE04goXaxWYtgpWj39rwp
tRmeCf//tWpD8tpJshek4sw72fUFlumQ1Jg3Q73I8mE9lGewoQC7TBM7eDiDxIZ6grOAxO62saRe
cfzkjfXrMuPFjWtf21erXWNkU7IM9KTg1NGDIb0AwrPzTiHRwlIb1O8xyOMcjmp03RVSlu0of4VE
oeTO2RPbqQbvi90id9vjkk0lcjD/DJDxw+f6GnXCevvppT5DfDNclxyJlEVpKcKbTleK9cRETqnB
eW5ZhBCdZcQZKpTNwA9dVV/mzcJ0rhFwBc5hwTV7Ya9mWKSPD+UTTo7Y5ir5u2C8UzbnYpsBSlNu
C73yLPODCwmuScVAJePw6/eK/vttSec68trA+CZiYGbFE5jP3hX4y5kDRzsR1spYlrEVQmhUfZZv
MI29YDCow+id+2dziGnOEzuV8gC/b1Sb0fe2f9mrSvJNPZsFFsHXmoEbctIUWMLeIu7OC1qMnT8T
Ql5yfWlYIxmpla3GBfOF9mJzEUZg/3sZ2j4GsZvNbyIq/FVx4O+pveYQ5uap3otQlh+o9YzlB/Il
hSMYF4koUYgVw0iGgHa2FLFZ56m1e0EOhjOMqEni27/2HJT0wPw6dOoow3oFrLcpEsQQ2fRshRff
aEdG4SxJCIELx8XOcstAoxaHarLoVwiS3a5x/8rQ7/J+3F9ZHJeQzgL0Ijf2egPeC4G7vqxw0ZOL
+AdlzngFKgFx1DzVAuBAc094/zN3SkK5j+f7jNXgzK0zjw2xc2Pntvevca/Iw72S50l+KVZH5R7E
ML/aTHm0yvl0u6oZkwcbNo+L9aKgxKAxwzK/O8BsjzERmHTcpJHv/IqjmWB6SbgoqEUZilFxO2X4
r7eitxQNEouWS2zXo82dusRMrMolmychaQaVwWIIlN4ZTPAzvNTMvYHjXcLpj/hRW0kZ1ZLOCXjG
3pe+5LzVNsDiM/1m5oWSX5ciOCiXBxlpfyMafi2EeXnwotNI3YJi7crPB5+AMDAI80t6IWf3x3d6
QnlitkrjeS2Xe6yxoKLfq4ALGhCCmjB01lqHjFhu2YrfqnhhrLAURRlJO1yXJEW6zCIFmEqhDxKF
jG++5F2K4Ipy+570xSm9WJh/B4XQYbWULfxpBJ8t5zPTNcGpZ4iLoDsnp+T1weOshjfGcAd/B97P
kiM2fwNjJ9xmRgQrKDQJqjOsr+GfhohApzgGMlx/SJozClTbG4TztmzkXjIg3cpjf2cCcMOR0DBh
7irYCw+bchoJG+A+3o3oq953pZzsjFvix844fHEbve7aOP3+ZzZsxvac8r/G/25A/SFpY7hUXaUe
/DFCDbYAD5xNM8uPhia1cIVdijL1qmE6VMP2lSpPE5oiedFsJfK+kq+JOm+bCsM9kbJH5T3DNlrI
+aHLOkD8pEOB8/GxTjBGsl2rVVSpS6XvDbbRLStuQcTYzSsX1L+qbpFLdYiB/glO3dgSE4b+YEAZ
tVX5eoN495wZp4GFLcJIyKWY9TzAJtWmz6nMClK1WKY5fBh0eiqdEq7vm37+fd2sUqO4W+wwaMJa
XvEKPIZQYKLSdAjnrvllaLD/PP2D3c/8P5sRBCyGkm7ZXnO/QSjW+Vm8TMjgutQ7yaQ9HJl+vaAK
dxTKG58Ekua/BU7pk6Dfr3aZunKg4gdV/V5xEyobhf6PtgMfEtWdrnbeIVZekbgklqb2jqCDFDaf
GDb5U2R7yWunX38BF3CI+9Zlr2+Y2buUe1plWAM/W7l2oiB7Y/zRX2jb9zDwa5+M9OevkxIxLd8T
9m8TNlzN8g22DqXnLKX3XKsqsMan6uabsddlNT1uaFajgDR4FHL4+65Y/8inaZd8mdvbHhHw7wKj
jCw7RGh+Eh7IwUXsQB1qCrT2SVFBITXWxyBQK2UCZpf3BslRpI7cjoC+L+eP+q/vrDfZqFmsYKu6
R6vymu5L0YI29ozgpSASUoeLKfRpH56kjDUkZP9DlVrQ9AY3jKbB/jnJPivpi3xayCdeqmgcZWkf
UnixvgYxmkTHcMgrjXj8yL55Jvv8mc/QOpHHjhD5Y+aK8Nqqumdp4OgRLT2RTiKG4I4gTkNbxof6
d3URUcyBQeRbAZOtq6Mp3Q3eRBNLXx2NhFuGDiu9UxQXLw7wf3QCVhyGuK0ydbQKFxbEPNuH4PCf
vE+2J29nim/wq9iKo/af0D03ocRMdJvw5ObpOK7uBkkZ6NYkSQV7LEygmAN0po2Dxe/8Ch4MnV6k
dAGapf6aVvTtRyC4KwJj5zz4obrWeMLoR+stc9/YIs7rJM/oadqbl5kSDod2sx+a7EOD5yCpeFVU
evmI4uF4p5tUc0fUzvWpshl2BbPEyTIoPgmgLd+UvisyM4ziPsa9ezt/vNhWrtHKHxsG6WnlEfHr
eHNaKTSRL2Ub72a2g5ujB4hvFr8SiBCgV2+pnDL5eNOkuq/BOrQJ27ow+Xf8RYocapK9Van7Dxb0
ETKSrdecA8NdbokdbqAZXYe7Xh6plOFj8Lz+/n9IZ8on17pD+w6q8an+hGaNfv1WPqUlusUAfhjJ
oSOF00vWC/VZ7nXDERp/ni82QSw+vS7J3qhDHmk6dzmLEbCZu8ftr3qvt86EiwcNf/fP2ERhLJ24
3Wrj5eJnfF6XftRK4GVLhmyEkmU5PwKj49NUlT1tC51Rq+WhuO/uRkqRcKLruUWHdiADK6f/7rZi
NCIkIvd8kReqhK6/Ook6ffMpEjgDvDXlwo9qelA/jE45dtXUr8x9pongCEcYUU/SNhWzTWoTUJkl
+84p5igGoOynjZ/XPx/KFtQ4Dd1TZAQrF0UL+EbJuJbaKow38c3Va1llBxvn21GsZxk27AckRr96
ldFYbA6rmh/cAs6Ol9N9ibtLDkSvV+Jlo4K23hXsjIRrTglkOJu0YGWlnXu/Xre1TQ+mgk/iXZc6
39g7iKRicUAFjqRQXHyKkR+REYrjkF7OLIPJJD1KzsfGSJ6lRyrUCB2tSTp0jW67bqbkO+6gHRAb
pWHU3QRDK/bohcf9oj85o1gVzIQKQM9ZH4UudBFMqKzj8coci9CtSKyL+tbL8TjKLVIjocpTFB/f
nc1jwnn/0sc/1NQ5EmZRL3VotubimQYzFIL0Wr8xhg8UDleYbYcnK99p+vfsY7221AVGcR+Ykhhd
pG05Ny7AzuBWZI/KfrPP24hXJUKCANuGZRT1NL0no+/jnYxAjzfhLuml4oOkgR34HSno+yYdy10c
rk7+O1BgNSJNlUABD2KOgCNUh1ld0BkaU47rPn+LZyrzLx8fFKg2e/YZYQULBEaDPjmQDtvjU91M
kjnM/Xl0LU8/oaez7W66RK+DYa2mQzT07JOJhzT3hgLbOYCPCVB0W2xcKigYkvhtCzsMMi7x5CLm
T5GEYoq06d0dbWLjSctpN/FAZAZBYLHnU9zIU2YYfzRb9ezmWLzyFsnmNm65wtYHnY+UW680S2VU
aUTA8Zu+It4ZLbuWd2rJpq69rdknauZE7hJGjtckqcfyvHeY5Hfb7IaACETLdny7AWVru3mF4ZX4
eXB4wUtnpOS0CuN5ZO4t2Cq7w3Fo+lWcbM4aOWKB65RNgsCh9IVbH9AxddBOry952xlM/dBSU+4Y
QJXDx9eWy9dYGv19XnGHnFeFkvxlQ5Xa3ImEN9mZp8/MbTeCrXTIGOpemf7ZNSd6YbM3nOblfeIg
PiRgh/54+0+ldWAOJZjOEIZ6hWMrljMKYubBpKudtRzETRZCI5sglrOoxz3kQMsnXGiVPeuJT/u2
2I4d+d9EczHnyaLq0lCKkPbcJ02B9ZgknHzBcfacVsZY+xzQuGJZx5IR/PqXc8y7lPkf+tUY8+4R
/kKBGetwq/7kGuzNvalU6PtmFwD2q4xVBRDNUHkJQo/jvaar/SNu+i5/k3WT45GRcRCGqW8AoCIT
eDOwTFtgHwzPPjs31gx6q7nx3IloVAz3JdradGuu664xgYh2/WZP+Bq/tJhCshpqRAM9tFbJ3O4t
tRqp4J6U4SRD6kW+vRdMR6voNhb4Q2MnpVjjvf0xVkhpFmeD+mNP7Qc405pQMyzjs9/YFBh9ON54
u4CQb84Gzywb4LyKz/9hrwmhfq/Tm+hhgYrXwZoeVWyMe80NVG8Tskt2BvxpBLYe1M1P+V6NZSk8
Trk+YkRcUp1XjcQl8VCbOfaZ85WeL0jvKuSKJjycwk1/0Ox3kh0F6kGx+TnjODCmZo4UOrTC3uTQ
7Cgp4VoYImOhr0UNhKabXknRga0/pZz1ovpU9t9TbGgk7PRvXVlX38U85+qSLCKcJImQBbY258G7
lSAEs64faplKZjkGdLmWh6b2TQL/KS8woVAeIfHqw79637De8clVzjSNcj5WGgdp9POFlLpyTAmY
oVakfutUIlyMdRSm4G5h491DJYvKET6aOiGpdCe+684qvmCzKM185yzO4G5HimtwcA0rJ4cEZYrs
AxOA7uCT+VUbbZ6vKS4wwv3qDwoYIFMxgZScc7peyb4PzWmylcRanHXvomxB2eu0ptdOoi5O3niU
ERSRUGOx9fp3Y9ZsScKPXS7K9onCUC7A5OjUEIbCcrcbiIjHd6+KWL15dBg3ubulUs9JyGsBTgDD
Gcqtrfglvu/RFWwfywzW+rFHBuM8qTfY33Drk1bRh8SF6iy5ZWxW2qRRCMbK1bL4ptkbDtQNk2cf
FjvLpZGgR2LPXobT8g4HhuO134h+wYXqvCjhbsZQ81GnyjmblFvtkedhGMPxrlSL1Bc/bwkgp1vX
a6gI3J7tSF9KBu2Revpsj/cMH54obdxGV2IYYP0Sz0MPVgEnJPunBGS5QNH/sF5m5fH6kyuY3jTz
pbxSARiQykM+bv6KV6kmECMg1MZ0B8VMuVeYHAjD9GMjXNVMsm/MKJA/2ouWdkLEGnIt5PwHidao
e+8NIvfTBJNPZmSYYPsE0EFEVajDgnNfK26+tsPcfSROtAFCwFYnA5Jl/0tDEeha3kdR+HRdQp0R
iLdl36Ikn4nVwFRKXrcjtwW4wuCnfAzfaMcx8RGk76PGmD9SoNQ4ZmvKMLgSbaa4BwxPkzj/+4mJ
WyIhX693PG88OL526H7lZka0PCWVnGRt+smxOKcLF7Kgpgqi2r5TD+UHj652gqn24oE+UW6LlyBA
fd0CYzqFyFVD7Lv6QXzq/uFG8ODbiTjE9Pv7QsK5TZ1dRnNg3q+9g6ECPoq76JD6RgYTdtH9Xs5I
dzqoGCXZCovEg5XC3PAjtF9Y+WOG0wLv1gOgbdcxMuRfxK8AKUyZW2gjpMjX9+oXLBQQs0Ko/AZs
Prx6TRcoHQzOt4uh9Rlc9DQg08Iec7j3D6d3XOt0Jk6Nhh360i2GugZ4C4BCA/2IWQEhS2u1sqCi
/hpT9S9JZv9eym6/1V/n5wkVgO7SlvPDhvCzd9UQAqiQ1btjm4GAnVbGjaMZgIdYwJY+JKKVWXD7
F1DhQzbzjQshrNIiOMSSPG7Et7OSbuVAKQe6k501GGZ1GBTmQd7UwxGo6ugyGCuJA+deHS9uARPy
A+3Tu1aDxEwqSU6el4XaY07dxJVvlmFBAL412FG5vXMWsdTeVym/2oWyIwBBtO1iD2TAEGeVLdTx
0GEyl65LNACzHOG7Xu+m7xfbkFKBheiusllO5c2Jx1W3CmRDPCc6rFOt4UB0B4KvGwuGxeUB24lZ
pn3cVAVR4X+q6K6NyTx2iyPTiXqs0iduBE4Laa65tf6JdZrwUBiVxz/hwL8VPUDkbWbxcu1+LRo5
AHtBu+7Gpst3mrkP/p+UQgtTkZ3JSgMxZ8ahbIyjzOUgJhWjIQKCXUvhAVObHiQdE+/XcPSTJY4s
LSpLZ2fFz2l4EXbexJQHn/FmXre3v4mLDwBx4xrz3iACg+2vWLloQazZ2IB6/LK7IWmtZj/uZqvj
5fj+kgyN0tuDSlTp0A2AKb24M/3EL0R04RRvd+MLloXw/V4X91V0ot2g/+7Sq6BWCpNK/rbfc5VV
CcEbdNg9hwXKrr9r/5iLB3nGUZrASKIi3jiBb2Q3V0D4oDpslPB9JQL3jMJjB8pt8wVcn3XCoVAm
Ob9KbRcdgaK1+elHe0SoOLyZZQejbz1ZDWXmRLIQBZ3MoVjNJreUjG/PTyKJMzbnVd9c/SW4YTJN
dFHu0GL9wivScOZk/pwgrttUksjMZn5tJt+GWxb6BN1MGVs1z9rNnArv5tkCW//iY/XtaPFZ85j7
HsyTP/cow6v5u1eocyP3G2OAAYrlu7eID4/pmNBUESMRexWk3R2ykyFfupzRNbw5Dv76kKz13AcJ
d/HCleM3K4qm52T8XhnnsAUXP95xERIQRq2OlKZtRal8X5fF45GJs7P62TNiAbYGON/3OLQEOfXD
sMnO1vhtc73BbLnEILfiGICCEbZ645B44uPvaPO6RdLrmy9WS6F8yQ4cTA6qWUeUu/Iu2z6jQYly
qwjXyEQk30vaKUz9OqTdCl5Lg4sI4WOgM8g0Xd4YQ8unyMA1LATnKU9DcRxoKDN9WC0LnE7XauFm
ZVNTAEwtw+weHRIJMjqHKrDnOpeU/ZhCN+/kqu9O5GSA9f3QWZHUz+DvJEcV6fWZjaqA1DWp3KSi
lCi/YO68wQOYrW5dpouTvbrWRPv8N1yW1s65MGICei9Xg4M0zmkMzrGEddiYY7jPBm6nyOdJ1vql
AiQKDHDuVsaBv4UR8KFHe88Uzytvfi5FjTc2xVimVhzSkV9cb8rWwi8HILJSywJlZi8BtsIKJQGl
y+wyXHPTWCmAzWNPmG3eb96r4uY2RBw1WTDOumoMUDPH1Po002p5CZf+KtTv1GM0e2A7zrsVE3N0
uPIafTLzOgpEjGtadXmJwry7xqonhfZ1Ig8HS3t9lZdltg3YPa5gl3pLMEDJR/KIO+Ze0RWrYBTZ
sQQwdeIL8poMnZxPAs456bDCi6HRryZsOROUPFJ2U6C6z/xFjdzQBQSldIDbGXorjWSN7rqr44tp
kTDfb3pcNNzrAzEd6XFMHUR5L8P2hFfwyEohlJCaSNEmGMr9ihkWlr/gMyhhUJqzRVvlIKGOhzGK
LMdq9h0VECYzE5rPgHVvkDAgAFWoo8iFoYvw5CW4vonfjFzB3StZEQlDVNfnSHucKy/2rqdBLoB4
Sp5O78HI+ua3aa1TqsQshwibJDG8NdRjQhbdSqNiZiNMcl+vlxwNE9srOLmCkSuSiBAFgDXjKkMs
lh06UAqNchBEyMGdJzfYLTaMZ74YRhJWjpRL1tCTWYHMtYs2TDJizv3vckP/C2XxrodprveVm5L9
SwkYmfeUPOBa4oTuaQCoobLAJhQ3PSlW7pAW5GgLJiRHEkQ+rAT+W8G4FHCqOd8/454Eh1w6z/ea
wv2KytPhWuckUGodGHxjC5g93UuvXFo7BqsED/aap9YMvrdkbpu/bPB8ockf+GQ2x2ENoT3+IlFT
fwzi93SpiH9gZHNSjmFjr4BTUEZS83v0uGUwyn4SJMRqWahlQcHPRfvmdz7Tn+a6spH/9eLZM/xq
py5WyadoYzkeBa+Hyz6g0eKv2Let7gAGbkBmXHOYJ+RdAbOUj8C4FzJ3xGQHf2LV7GtKbGp9sdjV
oUKgf3an1Tgo5wf06+cW1+hSAATBqglTlycJatn6ZrW/eamHkv2gYzWR/K6i+GzIjW9Piu4g5Em4
D2TuCx8D0zDR7bkE0KSwgV3Rf0q2kAdUPOpIHkovHbN9s7ZhsN7RDvqnKRnxHFzo9uXCK/sfekRa
5MXP9HtDmmHaS0yH7L0ZZxgcj2JqFeqwEzsQOiD7wR77rfkYCe4iRgcDqVgg9hdkXIdJ4ktJqr2v
dkHRS9uySt75YGHHWQAJo5IAYLXomsUaHj5cMdB0hti1WfkZXhMI7rlF32H7ZIZ51jzbcxb5qwMk
PWsqjHE7fEaFKp+47UUo2nupBlUT9DkZT/nWsRU7hJm1eFsPAFdyqe4rJnqudTLNVBTqgn6/oPGK
HnTiT3CKkCgKVMAqFyJpEvOQHA7ncadx3Jy/X/PodUO0Q9uX6sKeNFAfMbuxW5Qfdr2r6zp6Ofcv
qJq3BP9IhnNLEWP4U5n4eDFhC0eb6NH9TpbTIHmRlNo2HqaPOnV3FcjCF/KMYqJ7UVgYNCiKeswm
XEwuHKxbn3MxU1uqwDqY091R32ZthPiD+O4qvBfK/fidWPpp7zcMeZQ0G9BNCd75+DcOU42sRgtK
weoBaPVjOKqbcRTlQrpvgcBSljvg4tpyWYzvcw1Yz8kXYBqhIovYXZ6fbfwqF3piFvtBbeO5llmg
Tr+1FYA3je+YU4Mbo/IivJyKDY1CYS8C3RbnoH/D1iPQuUcsLq3PsdwHIVUzW8d4BpTxTqfgwUmV
6F+uNwvX1OzC/2UChmPpTt17TWqShe+X0oKw8HXMhLG5LQKXNaZ9D5gMLse43ktbxv9TDl5NRy7J
ZE2M2TnCLENMkr6VxDiSTifIBouxcSsClWpx4ybvaC0Bn+c291WsQdOLWM4OO3NXVWQ+leM/zjh+
3nkqN9vO853L95dRvFuCyYHX8pChIRWjwLb9uX9psjMuzHmjNnYOZUyOnC4eK17y4DcnR/gW3e5S
inO6OHUhNMlWjsWySz1+fTITPuLdzQ2bbIi3/YJxC1TlJNdEE+JSh85X0KBt+kKKcrOGsKHbjcnd
DhUVPDaAHNrj8lUknYZEltBrJzAuJThkZoLle0lapxEjwJEmPsb408GnBb8YEO4SwUwS8aRELGyq
NTOX3itwVnFMzb5a722wODPXFxmGeb096qy6T4VKzNYzbEDcrtLjDasRAThY/GSrIMjESO2gT9iX
MW29Il4G2TWtKTLnlx3zLTGXK/AmROJytma2WhaaEBYPwj1HtLHYQaUl0aRfe99ASXY/J/X9Vo4L
rWKQi2l1tphK4imdUVxhV0WxJMwKvEmvjNgknNA4Xda/cK4oxqN9/t3/wo2oswit249HY99tX3LV
BV7GJcLBUbvBlqVYs+rlrQKb2MV+vn2pUroO5ToZP5uC9Hocgy3d+9p4hwCAXatQuG5AYvCnUIuu
4ZaHU+BfeQtPFQUh6vZiYvnD/h1lpCg0kjOPizb4YEX1WzbHlVywdRl7jvnoY37BcCw6cQkBoVO5
K2CJ+Pkeq36YBLfiYfwhGUeU+M+YFw+cuVdEvju5Jfyglh6XCM4xkxqDiI9eqX1ys6d5SoFCz/z/
ySii+wkLN9o/feu23om/h2PVWI1IOf5FXDtuH0h0WymRyCuLJWh3NzYGa0XyYyiYuAd7bwdzOzef
MqXzTZ7iNFVw906MLtq9kmCL1fcRuI0fNFysXW1hYIeyU9MmGDam5bcd1E/hITWE+nmN6O9+Q/jz
CbOC5wUF8YszyBqrhCVEYKkn5f//D7Gt0LH6cUKufb8V92D+cCZw8H3vSrp0U36/o8mAKsX3m6yQ
sx74TTKVNYoM15lMbSasoW0Nm/4UDLUlqTQtjkGJaCiwrgKpMUqpGu7PMp8zznixhscYxd2WTBkF
zUctSUmusDpfIk20UnDTE5tjFZimjQqPzocRHN6cxAwLMnFS6TY6kB7cmGMHGHJv5g4q4ncUb6s0
JIzBCYtdt59ef4ta5K0CuXe9Gksz0R+y2omgjuXA/kqzzQHh5Ou6coCh0pDL976TaARnlxfBoIO5
F/RueE4L2Eo76kD0NGHhMBqMTmYSE5QuE/jRYus5GgIupHIjwQG7b6k8Vl/xHOR6uEkUBSGyi33b
TBswmVlTwlRuUMxyuzzd4MbFECB99kfSYz3yteu2v375VFBLQvhGVhnUa5+2dFpGUeYNyhISCXUu
oQdcCneS9jDy3AAVMZcB9T3b9kdxjqsO1iT1eyKj/6+hRvozceAnFREVcpkeRU4+WGG0gjyCeirR
EbcftJ8UTqwAc7AM+uVqQmkg18Hn216vOcnDN1tGJTjV8nM8wi8WbHnZRfXt/NewHVNDTaE7733a
i3Zmlnp+Td4ZoD/spWXBx061cD6/HAklw11paR8clSTmOzaOBRfUgvo6LwLFE3hTdS0uvzCjUFCv
OG4FTZFs74QxK3bXNw2Laz0OnpTND4SNGy8h83wCKGuwCZQ80HeZ4b5roxp0QF6l0A8X3Zo7SQ5L
jatYOdHSjbjNAej9WGV5Vpoljm7OJ3+E7HOb0nhdQVFKhOlGhC6U5w+c3l4tqA/5nJdKNAusZI2Q
RKKa3yq5735lUXlJnygDx7Du3YHYjsOCz1TfIImmH4vOpC+Olt2mi7hIq5IkG5WCg6aS5S3eEAJO
8Auj/Hvc7KmwfQNhjcByb5z/dpa5+mx4qaR/gNr1t/cX6Ez970fqcL6r1ehV41l4Tm28m4joofs/
2lKSmGrvnPrE7Lf6/KDA+C2rmfMQHMJT++QkJuBrftzgKVR1SYFRJXFR2iaC50RnN9iyXBVi0c12
guUYjMdQJyGmFVU9Q29nngePUHJXjNZ/3QoSq1MMSn0ss5I0FEfwD7avYwLjsUIfjRn1K43tSTmd
pUEe9ajIzk3H5CFPeUae2FDbxaX1BebhDyRxlhtpp/0UV0nVAkuj6jT5AvYJU3P512y/bB2u62FC
eS0yc8kMyeWxao1N9oq95Zvr3umrEd5yFtaBOnimDPvWqAR1nbWLXQci4nJEAYmx7eNVs+3Hq/UR
adKJRD68R8TRVAzfRK5qgrJ4Rh4412feh18YLhcpzd4sqjmY8aJkQ1lbrQ9KM2f/AeluqYnJU9AC
PdcBsBopTz5K+xliQQWfmlfDiyYLLEpG5whh73ivLJlb54AHFN6v3zZXZk4yRlRYwawL/ltga5vI
qI4E4nSdXO79VIUh+PBKaScoDVxqP4mkyR7OjGvlMsvpjYGJ32HP0f+XmQBXl0N/DJcMsuUrQP0Q
r0N0e56ZLF0BfSJqHlqtWWChTzjcoSsN5ff0RQN/IFybxnr/pnkKnTyvZrzuP3IAOW7LYJLcidqi
DT+22UZQII+n3hkByh+kFhaHGtBRLvNjGDHNcZUtYyy5bFXprsByHE7jwIFK4OdIHfeQz8MfRgMv
ngPhqswH6rJ0yHn1Aj903eJqqHYW2f9D5hcYKy3ORtooHQje00degx9W/HI0oqgqbbtX69InGCMl
mO2jRE+q0+jHID5uTXN5lHSuRKjAnFX/v6EX/dlFLjzrKa0mJmlwg4NNlOx82jjt1RKrzNQMyM29
FdLRaLmNeADVfx+miMTq9n8MPOVf/f1ZKqOCfzLOxYmo4IgTK5pJ1DbGZpiCSlMaTXBo9+PPlv2e
qOQu8YB8c5RM9BoheP3yLUqQphAc5040d5Tm8W+AGN7/4tubP9ymfW+s6WymAQvZ5Z/+f7TLPO/l
B5aTevaFkwA+tt/3YJuotWLzPEL/Pk7xpezlpngkpvhEvpSGkMXEKoxQVDmns2Qcj9DFBhThwtBf
LpPdjbXe9y2/K0N4i54FRh5QAeyCGoZo43mVHjQf5TCG1njCCSWSdq+nPBVCM6EVr58O2+yPL8fv
QX30/JQtZRmERjguqwZAOkzTNBtnzNKoc1PvAp/zW7ecfWgNSAtJPWzvtyxFv5BZBy0i/fLuXD0/
MBzmQIVw3nGLlqWxRVqlb0VJFY85fMk+TH9+4Oy4Z0cWwZ8m/6znfeLn/ovRj6WR+C4Sn9N8oIyf
5Rk+ydi8jW4AULnWMrTyUGEXEZD48IyYPN+PoL1t5cUgjuloYzRLGnDeVfkZ64BmF39LQonHjDae
jHyc48aphnV3EzXGNVV8m3a3W0PsYCWV+i+L/KkppxYPktuAyyciGR6L60g7GQbWouy1pt8Xg4mF
d1fTuYyNIBUgEE+aK+GW/cBi6QzFm+Y43MCEvgYA1ioqJ5dTQ1cDSQpNR9D/aiBgw7nINw6NjXtO
9gahP9qL7h8kYf0NJ0sEdBwnM/4MDVtwdy/5ozxtVrWNwt9XTQ2MG4TzqDQcHuoS7ibctLn3psNE
epxWYSthRK6ZgxomsMGQoq7xKEgSrTTwciQsK7UtOeowXZhW5Qc/2Y+5SL7hScwjdpD35YkcXo+o
8RC0Wa/Q2gdSUgXV5ymWbliCT3iUG7VIAhu1oGSU+8YnUECLdZ3NqiVUX1u+YjDrJgqpGX9Kgo28
50AWqkLkLv9Or0U5EdJBGcu/19Ty4QzAaR0NxYH2TF1ASWTGu78e7Abo6pWLvGehxOFqbbKkPm3Y
8opRuDKsxOuqgPsw8sr1XrsGXI1wsSiztkVtdAe4WmmaMvzInRYXQEd/C+dkywMpBuNMKLD8n8LH
7eAIYrjpA1I1ch8g0JVE73g4H7X/ysqBMDNeGu2SGTmaHt46cp/IlwJvsbpNGmgUKmlsdnK0CDsr
5a1y0PJO4j/mUIPJyH7DTbD49wD4sSIVN3vZSVSszGw9TbmxdC+lwwSPqQeWJCYLFYvBQbwmp5yo
MCJsW0tgFBOfrAD4mdhkITTGjbAaUS9uNKwZBiJeHgvdRBgua6ER452vGb4GqbelA2E1MX/GzMdN
kYSG88w76G9Z/pmVTm0uprGbDTQuGUuSXbStk4d+y4pJ8ff4kpKwbE2/zgFP5A976LMBVWGjdZAd
8z0BCOJ1WK/Z4/0Fxe7j1XFUlLzl9k6p/RnR9OA9FZHih2VM674MIPZkkdmiwEjZObdJGqVXaTNz
xchu9LCGHWIn+0tOKRqX6tK8rVTzL/MLCT4VeKUFcEdp0ps22HFO4RNnIB3+wzBZukrk7rIa6JyP
i5cTo5P2GnLbzdPFtHGFXAY/i0uYiEnMLel+/n+g5mUDZNBYDd5VtMWDD2UFZa2ik0IVSS45B72z
xswDZIZ1dTu4rw1h5MDC7lN0AvfFPHR0+GkpYqI+LlccvhoNToYiYRXxiHk4nvUO6nfKIVztpInR
5HAp6gLC1neUSIskavDadhOkfco9kYM4MMCt0VGsLENQyPjjaHzLtokFVbu7iliXo4jAR8uWH4qy
jFCa5XF/9sZvjgUZGt73DjX+8CJ4T+3KdioHy38E1OBgG4lrwegPHiTzHIGBmxB/VfZJzuYi9I5H
DzWDf9qDmPJmHHW+nfyHYL5xBeucG0spskFVIsTR9beHpRb760mja+NzQsT+AZL97/ACAX0SgbY2
pqBxK7iOUYCQ8t3avjmuvk1g/2hzjB+o7liqzSadupP92mPG7CH1bil9TiBV/1Mh0El9PBs7pSib
VfOSnuaZHbiGck3JqfmiGqHLzqXhi6eFseG6vogTQkt3zUhUTVQiJz/LMvn2MZEHLhFgz4yfD45z
p9ZHi2vLyvDYeAvEdchMJ3gBJYmMSadIp4LNt5Gt8EbFOZilKGBDmxhNhOvScu/WyP+3ZH7KV6Jp
EFPtsE310BbctZN77+YSiKDlP0KVRqOMJJV0UxH6iDfgkpJWNEGgS3PSNdrr/zk88AlrNRLx7CjW
3yDtx3o1MMGQfrqZ9N6xfc5e2BfsmruvYGtrq3aba1bonpylinbvvx2DMDI4g0rF8BirO5ezKojX
yW71V1OVBXJ3fJDr6ZQSU5gdI97uKPMshpClEYtoteqdcWiRChybDXkmSAsCeNC0z4wj80ZLRsPQ
o5eWWIm0LJus9TmUWtbAPCRx/KB5maMb6xFdHO7QLFRvxjflIfK4tXNv0/MD8jxMwBcJCBvZOhSc
xpdZVlcPmA0Tf9s9pbg8nrZzCOIUPvZBuTdDG5n7hwPXsiOYplGe3Fqf85InKk7TvcsD7etjMTq+
rD3IifsnfrpFKUANIfWTChHS6P6aPZA3TG6t8UxKDDqFXBfXpwvIm/Ak6f+Xf1MkDJfRIl/teXpr
2zKHdqLh4R8lUWjDHYB+VAecRwS1uARBZgSD/Y+d6thktrht98VAwNJY6c9tT2U2XvMBFl2fM0Ms
ybVd/5It7W75pBiktSuDfY0VHWlwk2tv35BfAdo7PtvFBmUssBjixKXzWyQS+Ppdu3ppxt0p9HeV
MQXJMeSczRTgr5blJqKstox6fW0NCy2JGmrV4XX4PHrqtMoKbyCayVugLV7pIp8eV9hpSgSCdFAq
0UVRcwyGyexmuugkvrt1kFENH05Q8SqHxArQGA4+9k6rzPSM1MDE0sYWhJf2M0IWRQq3WgUjQq/O
IlwXxHLPExVOvEMnP32lacmNk8OtEoptQqiqAne8KDZ25p5llN6plC3qPtz9gPfTX8s1Gc9I7Bdx
qRmCsFD47o5vFnl2AQpSr44CVS3HAGmqqjoqfsPS/75aHE9lE4lEY2S8kIfxEVQpFvN9p933azXl
+o2AuK2ks8U3yRMtNs68uhYqAjptWQtEPfg5lf1/wbUDx+K8JgqzR24sXee9MQ/K6wSAnuI1DkiB
5RXQH0ttGD8v2skCkTq9oyOwvl4k6Xdez4/jKw/4KAb25QZ9wnRb3DB2lmfvjmWijv56D3xvgeyP
fLmIg7c7wPVKWaER/rzYa4FzxoqWgbwsolKyH8OFsx4Q7FELcAn6jSWvHGmKRQwR2I61sv5F34J5
XsO4cUUMUIqi9H+aGZdL81K9FKp6qmg0fZsQAcHBjM5xuNHyOe6BzcNZvdzF2OEq85s0OHXL18E2
EdG0M6z5wzs8vUrCnS4HHSDGbLUUTt9qjDiyFthwklkGDvjQofzilt/X2MOjateegZ9kM+/SJF6E
kLpwR2mQM5KvM78lSdnX+ev/qh8sad5+TQjPOO+aQs/m6qlj5mwlua3aOopShkcFA8RLsX/dDJWQ
0jeejru3Zbb/zpVY4i/0h1BkFCaoEqAV17rLn96LNuRLNl4/Yjiaq/GNQ6f2kxD7xwVkZ7F/jAiZ
AEw4ZXzsFI7dhSY5OeTBbdje7yerXMT+k4aT6v/sDqdODM4NrYzXrPJdCq+dn1zgUxr0R+xyvkHC
fCR7+9fQpLjPFIGm+QPV+/ODO/GXoPVm2Q9RiehYSrWYangwjmG1lYqMkbWDhLP3cqSfhV499fZF
ggKNuHt+RgqR7USyt7cb2A+EfQ30bFsM3QwgHMHKBfWewKHqWTp84AI8h697DEueGNAKUcGSupLF
hfneNgoPkMrcvRTqoTLisxVl2PN0x0cKIr8Q49sYTf4ay5t8ig7UeE0IF7YJfS+2qHbK6FRYaDQo
+rhoQoTVoJQg5YQouGUSEJRnQG49kds7oj2e2MFZXk1JlaB8YJa0M1HRGSkux5FcidBDdNn8/m6Z
glF9+G/az69xFXS0ehJZUHfHPVt0Q8m/kitdoY8M7ZrEVluahBU0p6dvXzPK1LtZFKB4Pc0eWfmL
yYQ9KjM+RltQvm2UDOl9e5Lw2NlTS0Qhrd3njNKBemUdX2fcc/GfVogOHESKwMzpsSE+sNQyRcp4
usk6PQuxFzDaq9YDxPDyJODOV8IS1gCRRRhXM1ohbs5+XGJjrqixQ3LUTFxnCh0WLQ6Xp+BETIEH
dt/fS+RloHvCx3F/e99lVw1bbnZxUBLGhmOdgGuXWlVfNfzZtewTPUuTxPuM+6mS30gwEyes9n+m
0WGQKLzzqHzYFlRPIOHm0WhXYWZ/vQhZ6S4U5Jb4+seoD9WJf54x5OOT6k7U+LZJvtbcAhOLRO+0
zzX563QT6WpmxXPWQU+TMpAQ4W7DGgIYXKdUzDoBkaxbI3aSeREDSyJMe7IKUYxV4/fztgKjRJ6S
X6OgC4krpsAXpFAQyHQ5chtVkZNKuLP9idMVH1O5gFck+4oxypk9S2Lz+vbn1d1RhlN+8+WsNbuc
a3eNrZLBi8IR59u14LL8rtELOEo6Qn+0Fj26mHin6D3+6L/Vg7hkqoz1IBSEhqyS1jLsDcaCCr+S
PlMTbKvDRBaN0F8/RFkz6cjgP57aDfk50EfmXTllQPxvn9Ju/tiy16SgqkzSFJiepWQ7xBHfgulB
QndD1+sjyLdTpMJEOvoxtE1cZ7cXEpTZxjjpo2l2/WLKfgR9BcClEBrfC8iqTIGwQfQw8x+/B214
UXKp212LGcqmPnDuxZeqgCAndiEEs9fLIYBZqurtiVOYJTJ7Jb2E7mXasgXLCoRbMEp6Qj7RwKqD
WKVESknmgW7uVgR/MTo5azxRREKcWu1SQtIJJaqZNuPtqAcHH2iQ318W/qRu5tMaocgGegM8Okxn
vGnKX5963SKkN6+hvNMGNCN+RsxYfRSeNTCW0RrSf/aXsnT8YzjFEK8uVJs8Vkl9t63q5ksXVp6J
TD2zdva0fDRBH4o0Y7IisLF7g8XuHJR5d/27Ja/KHk6fRdoK6QhOI1ouCyARguDj2XaVhbWD/7rL
CH9XCdFFhceFScYxEe9mxwM3dRuSCq9dKmJBshz9Z9qnCq7X8jPBEovbaDIbNGj/iqx0cfoGeXdq
B2TDyWTyLt8sMUJslvdMXytFt3XyWX/5POtQAFgrCu/HhLZPnriMBBmkzq6eN8RAJtDXGH4fkXbG
piPI6cEqwVrZub4InlxQMOT6svB4UM7ycqB5lfbRQ+sPK7czwBxoUXnQYTnGMqNRJpdaJvzNLIZl
8XoK7V6jmfwyccG88jcTXQk4d8OzoEeDuEo5Lpyyq9UWbCFyAcpA3d7TNHDNvrUNuPv6YkgAlYYN
8F287O7T1uItbQjLNvfBPGBZt5V3oJF/4LHhUBDYhzQE7V8YfZ8oMzMMGj6+crQW5Iik0K/CHry8
86kNjiQlU4pHzAKw0nZMj2eVuFFSSNlpU44rYpJ21JRQ943ZwA1vVv6oxM8zS/MEAk6WF89dPtHj
dRNuiCjcF7zBFHJoHz9o8O8P79Yp2OBpcld4oVeTOxPTr8MWaQEeLFkDqlas7zuWYktA3eu81Z1F
qRuu/g9n75JbvqVaHX/e27M/kbQT/iioXGL/AzM3GARnyA/594fPYW3FGqziUPHVl5vOYCBg8KP6
269xFp4+1tQUEDAXXHnbpAYNj8x5FOSsCrcT92q7Xnxcz2OblW5b+fuWmS/ohkk+eC4I3YOz/HRn
uNBALS0F3gMdMZjtfvyfrdeeXI2gR25eh6OzOxIZ4Z3PC54sYu4vlEiUJCnmcyuR1VK7uvTI11LJ
TCpcVT8JDiURJFyI2H7zFk1pBlZx3b2RpFWLFXomRxHCPhcIabFuknHlU1WxYfli8HcUbgc7Q1EY
cWR/0/MlZi67pk8+0vlrY0UCba1VRCWAu/I86J+/4cmqT+v0fnHlYIV4JvvIA7kGGr/Ry0sq6Gvn
XevKmA+Ld1379Ebk7NQCprXjhqcB/4v9KQsmuScDqoO9jSZTxobr04r1yeEAsHeumZDpwjmZtqlP
IgXxe4Fpwdn9B/ZNPgcKWsDzreHkPN11q1HEeRTlN1KAoAu1Syf0UMbFUZlWH09Ssf0p/RIuKL6l
iSWrV3BCMXH8y1/4gxONmInafDPX6n1rEJ7BD/1aT/7jqptM0grohAqOtNKYLWws7fYkmWwADK/R
jogPvC4+JKlO25UlQSacNEZ8RhhdI3azcwGXuHbU6YEjCT3CETrsAvCaErv8+XP6OOJWQjkgpnBY
gdR84E3uACERwkMHL0BU76MBn2BxiVCUeEVkMR+WVQPJbiUB/NvUD/L7+gEANMnGRKQ/h/lNivZ+
jEj/8l3o+3PRLnJRa1y7Y6gvtgUDfjlRyO2CJO0ukGoj4VyoUlWD8bQkkkO7wGulfnraTIJQnMft
ml4x9clfexUHoA2OK59YmzcB6wk5s246s+UkrupDuQpY+Gn+CgU5tf2EOHMZ2e41OMDJ2SrSsese
9GirHaj/WW4KWIuK9A7Ye1tfEEpmMVhjW36oVr8pX1faTbO9MQFtlnhP1Pw3lf5AEeN49yjE/g44
VPQVLKe/Sy49leL5u88miXbkq4j4IgucYBVKrfx59Ijpfjp87cc6DCvVU9Day3fFVe6DN01EeNTK
B3Tca6BeYw/GD9pXx91nU1iWGHJFJ4QseJJXJEmFnMDP/YLX7nw+5Ql4tV9CqV7U7kqCHqb10AeI
NONrBi3aAgQ069MD/rba6am68gJy3DYwm/mPTUsOGDeExw90acQGt6GC9St24uJNUeUpvhZrZyJE
6hXprwISQ54CTH1UrVwYJaLErm3XYHf/O06P4hlIIVxnBdNl0RjQUzkoMJbeUJ/bZY9LkEzrn5An
txs0Pnh6+/D7ajFDfjIvxMM5osG3DTgTrfFqqwMW7Pc9Yj246yRF22KWS7AVoMy8Nxb4Op8Xu2Mo
pM+L0rRJ37ydAKnMFWdSCoQ1aKHW1a4tHnhaog4cSqZfXLXzyuZBZcDH9i7mf/A+hxltQEyNpZ/F
bQRQN+56T+ahrne+nk3W2ovjSbL9npl53v26lU6leMd7SZDKuKMCVUKZXIyisaT+ma3YoxUpLP/s
NGgr+suCjoZSP2UqZtaOdSj/OkPBK4vsb3fakqMgIGQKSKlvAhezsUQeJK5WY6G2VVev2pKyY1Di
q6rM6aeFnnj1HydYFXhvtnDSC5p7186i0zFPLOtUfIsyhPfOWI/Vdlf5Ah6/TLZsNU0ELkV1RNdf
eh3ay2Gumh6Bk6jMDLGGiCCdoX6U8nnL8zqfldkm7m167SBgmbtgrIc/gmAObTQyFRtxEdRPdWkq
loUaOrjzYUAHwr7LUYnvK0jM9LzCDwx7qy452mneQ6q2lw+L3J3C6c4TfNgvzKy12ij84B+jstNC
pzK3f68gB9ElR6q7ec8WlLvMmJmz+qJY4xRS/SieHdxOpbXmTLN18SSufRebjv93DcOg76xeW5mv
3W1o4UifhIm30aUsz4YmLum39TnoOnuJrXXeGIazygeE4noARGA/VsknTwKxZ3R9lVQpPZVZqEmG
WTj+Vz+0eaUNLjUvWfQl0N/BkcOq1I5djsntksVejdBoerEmZ19jKBUeBNPkgb9b6uJelkxVbBf3
6w8UHSH5eXD9GWM+S7mxYeiuC/onBWtxbN+EAfXbIhfieIbb4s6bB/aoXZKmsM7iO13/YaNBLFKC
9dwz8tu0KiVCwWlLxRpDQnzSOWiO4xCDXRQRXZyl3z0HUkgvmr/sOYt2bh/2KKslr5aiFZX9CqkR
e3dmwgnwnUlWyE3D0ndeRXRuMbn7UCNYoRZuNV6Q8FbL53AP3A4xV7D3KLdqrLDVpvWbNuhexgeR
6bLe4rRPjKR3KQNW5xS0rKLFjZC3VPgm2uG0Vpw2Wx03jJdk/sXuhntbDLCAVExczR+jnCWSGajw
aa5vcbMfK07k51GUebnaAEuvCutLItwQjpmRrMqiTJ2qgxwKmI2s5O4pFug0+SWXQf5tX3YzrvBK
U1nbChyIHdQJ3T4FrqtG9qsZAOfiDYR6T2Vh9IJ4XtoeqHbx4nfSSQVYRP117cbgdRlAxmy5x++O
YJg7KDM8F95/GEBr6f2+D/1os07mUNZ5i+u1gxfUVCbCq60F0Zr5/mBLchR1qv6EeMmlML3s5tpa
5rEvBbdRebEemDmRNHJcyuToXI7DkkAJH7SnzcIvjdxrpnXFnYdvk31WYFaOHCxxihUQzrgPjXwv
q0B0Yuzv16TqsElKrqjtrybw9L89JATlTdnYFXjbyxHujBpTwotjpmuI3qIQpf0IKaJ+4/+BzHlW
z/4N2iSNJ65Ojgcvlei6c/rcIuS4T24go2xwvEFEs9Nsb7qEkwvSd2noWSG8FGbuGAUmxBAbnlsI
Uy253hWjYTRmJZoGlBoT/+PpzMDJglmUzIGCOlKA+CteBLPuJziOoOXCovHjhdfjLhvO3zdMx1hp
R46PQGwvn+uDKi0ZtlhBfMHkMr0NdgdEc2V1vEv70e2Q6UEJt7Gl+4EhgCQJju4lDgWTP+5p3kna
X7x5nSnVtlhmwLCtqZgVL8+1wKTlgtuIi7XZq1WJ9C5Eih24FfFgcxtI3WKPW8UfiL2P31npkSts
DCqHWrPWq9XnVvaRx6KRVKxtGHThXcE2zoii//rRu31lpUva2kAmCiyw42XkvTZbyHQ2YdVH/gTi
puqMCp/uHr1yWpkkSn4NeffdMs+xqXbwSDKxY+P41V+onPrEnebRXn1yUHfc7lROSTquhk+nPPM/
hQe1oBB+QU25HRY7rvP4Z0b+SsqC1SgipfH8cuqATjHTBxz8eDatLa8OrxyedfJmApx+tMgs847B
s7NVSnVLJG7guPZMFmveOqTr/+Cpm9Azy0sq6xDOEGW7Yl4fE3sIT8+mbrdLsSDt7FcPhy51GObp
0FUspYIxGuIXKefNCqPyTI2n1s58JzHwIw3GQ8Ywk5lXhhnPlUeZXjQsbNhjNXtppvVigi0Y40Kh
EbrSK4EXwWICnW5tO0cQf61Re83cRTJs4HU+JOywYbJzvBqhDs/B1AItOUNui7DcNYAICQd+egXp
mDQT0u0i5EavoXyfUM74/XzKZr5Uy0JQIPJTh5THBxnaK+tu6ZJjqzN1wWjun7Y9TxkaKQO05rtD
wk1S+xFjcrXJNJMGXVTLCGHSaZRnyxP6/6euqiMi/ZK9aCRaoDkrwx93aSSdSg3HWC/yWH1VL88E
CjesebgOMGtgewBnFvcE6FG0IGrHz8B6kKrlwGrP5XLP4mf8+470ZEWM7ttX3nDFuUQTz3DIdQif
KyOEVOa5w7sPWoIXNgzO51CqZt5awROB9TcRD/2qtu1PXLPcfuG8ptkGWrxKoZwyPS2PlbgsBMBv
eVSgYdKefKQqCF8vpmWTE1PUauxJuUbZw0NjvSjlaYLB53cyL+fkxatqezal3J424iZM9VkeN+mz
G9lSrBmyF2A0dBwiQcbZaS9nEvTmtc6ppK2oILvNMT+vLSsR79nUrJnKAKYG5Ef8a63xpdmoUWoU
DzSz+vu9mR7MZpLInXFL6aP0LfqFfdEaFxH2eufxB5nkixWimPSLvFqTUWuqwmFHwZZlq582EF4V
y5cwVX0UPvgFrDPm9U93EY4v3YNzAZ1DzIvdiPGbGPsSytx9PU9zggCCiHNx3PJuV26Irdqfkofb
SUODOLZ4vSP/yBisR4RNkG5eQTSYVWh3lQT0dmVgFMWze+WxBrOdh8245m55vkbJ1mLNVXkEMjAk
cqERZGnaiIvoQYKd5wRChTgxJ5cYseTaG63sE21ZPD6KemzcEPNhA7O7PUfuQKo6c2clXaL0aEAd
FMgexNFTkF5m30/HjZwudREPP9ElaDKfXBR3Stn0qkeQjNuA9NLXZkChu2tV34epsuR07w57GdJc
nH8MSLhDtIcmAy2FDUTMkgfvSzVkxeNyk92UBvEqZW25SYlv6cCOvuvDX+K12NM33dWYsJZGO1MK
2Sq2c1ld+oNfF6g/0zVrAh7jpJ5G339rD49gKr3ngis/3dvMAdufeP33RbJwwl0CiPUY9cdzuIxb
zcQB7TyrMthHzpRe4AP8o+HV38Ios3ElNr6sd9C9mIKGpZlvsgN6gdXbZjPvPLI1NbF6tK136St+
1eptbJxZbZWsFuh9kN9FV49SdHYcmUOwSRpUKndQa6YIaFCzH5TjqagxTYMMVb7rf9h13K0TDk+p
Qsfu0IYSSGECYMp/U0HBoOaRdTQIMq/eQnpv31//ohT1oAf2Zgzfl2apfUicEYgm6Ok/qW/RZpZT
6g/nd+ZjuSd9b69OKjV0SPxJ5To+8TtM6GZir+wjriXskh3GcYNx3rP+a7HvieiO+8ZCsHHMjNYx
2SCU1fw/sjQ4x7CjOROPx8/Cw+9pKXfY4Fy8rGCmGQ4okir7x61Gz3y9PEmv0PUqZQpchL37vBoQ
3TgniBwUThmxRJaTTFDKxU2+yhgFudF1+rY2xISZX7ewUO2fF/NIL70Awgs0/aUM3uEH6jp5ENa8
rPedRFbUTHfOGD0FuewzNjtELABFm/HujPfgIAxXqD8icOHpuFB/urASsdmq9KAxynITBzSkUzS2
BmxSAKT8Y0EF0sKxMTyTdhqi5LhRlKW/0N107Eba3LAUc3qhf7XlLy3F9D9w800+TDxmjt2KApgu
lSzaZt8GCgKr+n7ZXQb5skals4baF/mJq0G6NSXGJganMhDOGmfU4WNLmXcsimokQGaz6XQn8luU
DfqN20n68hOAZwChWPEKn4s2UXPZzA07LuSOuRsxkZWx0H9eZgKrBkZIXFqADcdDN7WCDjDe8cBw
oC5i+j7p/scQ+jJwHQ9xyrAuBzYmkqoWYmcCr8anFJz9/3XB+Wxl85GT6z9JRAbq7mqnenoKv2nw
hZOHJ1E4kDpJC9nHaJuFaBtclA7h3O1v/KHaiJN/H6x2wmqDbN+yvYd4+b6X+9hjSuu5UxmrGp0x
jmtbH6rlMEd5naszUxzn8jcjAs1MeQ8vHr6eDKtsFc/iaupd6vJbtwY85BB9sBeG/ILItFRaR40j
xVEaLQTXe2GHP5hkdEOnVoLJimjRU2NxIGrEM6J6MKHihhMyKx2wxorbVO6+y9qSZn6dRbAENd1R
LDS46wJ63tMaw58UJcQ4fx1RRKmTIALhlYnx44BYi7v6hD5pGefcXoFrFLWvizRypER1d2PDcoBj
nkNOJGR8LgbyOyXK1ukZ+ekFOyiA0KMnlKuFSuPxgk4J3gyX7y6GNm3e29LQl6gSt3pnCmCtVQ+I
7ADHcTkzhEE2B8IDQngaSOA9llfV9dJUnflekt7BVQ8KJAUkwNlPa4aQ9lM00NutBRJCXS9zdsk0
tHvTbiHc9a7ixahTrLRYP0+FN59eif4v+jzFesCL+OCHWq/2krz+rJsXo9izokkIiQKGH3+Ku5hr
o57RpLI4ZRNKHtR4MINgAHFvkrW9k+IvP/KhyxTgZ6CvNEJSkPsrq7J5owhevohZUeUH1/4+gMJB
YpqS4NDihAXwCb5mLZz9UR/4KXXDR4l315r41PS1vzBb9IcwU/nb3sK5/camZtL6WZSYOST+I+Dd
Y2OokyosjKnY7kEXPZb2kAUUIE23VP6pJZYzvz6F8xj3O0If1yeU/wAcEqVcvnAXLzjO4hCaUFFs
d2uNereuKfPjjYxW16ZwIQ4f40sw1rq8hrmSuPK3692iahbC+VmbP/mnzxfdcPkKajWSV5Hw4cFg
rsu3CWvTpY/pi413lnDHu5pNuRraLf9bRHqllkwNUg/AW4Vl5h7zQym9NOXWNYvcALabJakuw2jT
eXkqTRfZyTl3XMYf7NDs4E5aiISOn4JWhsnTDcYMFx8JpVlfEI21TqWIRpASMqoh2smI1RP+6fiQ
JQtQRZQ2XyrogtkYfiU2WpbqcCaDh2dt5VVR9jwpJKKeg/idYOlqvZbATSN4PkQCcQzn0onKUTM0
GkoxVF/IRbgVA/GdHjzR0A==
`protect end_protected
